// ****************************************************************************/
// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// Description: 
//
// SVN Revision Information:
// SVN $Revision: $
// SVN $Date: $
//
// Resolved SARs
// SAR      Date     Who   Description
//
// Notes:
//
// ****************************************************************************/
`define RANDOMIZE
`timescale 1ns/10ps
module CORERISCV_AXI4_ROCKET_TILE(
  input   clk,
  input   reset,
  input   io_cached_0_acquire_ready,
  output  io_cached_0_acquire_valid,
  output [25:0] io_cached_0_acquire_bits_addr_block,
  output  io_cached_0_acquire_bits_client_xact_id,
  output [2:0] io_cached_0_acquire_bits_addr_beat,
  output  io_cached_0_acquire_bits_is_builtin_type,
  output [2:0] io_cached_0_acquire_bits_a_type,
  output [11:0] io_cached_0_acquire_bits_union,
  output [63:0] io_cached_0_acquire_bits_data,
  output  io_cached_0_probe_ready,
  input   io_cached_0_probe_valid,
  input  [25:0] io_cached_0_probe_bits_addr_block,
  input  [1:0] io_cached_0_probe_bits_p_type,
  input   io_cached_0_release_ready,
  output  io_cached_0_release_valid,
  output [2:0] io_cached_0_release_bits_addr_beat,
  output [25:0] io_cached_0_release_bits_addr_block,
  output  io_cached_0_release_bits_client_xact_id,
  output  io_cached_0_release_bits_voluntary,
  output [2:0] io_cached_0_release_bits_r_type,
  output [63:0] io_cached_0_release_bits_data,
  output  io_cached_0_grant_ready,
  input   io_cached_0_grant_valid,
  input  [2:0] io_cached_0_grant_bits_addr_beat,
  input   io_cached_0_grant_bits_client_xact_id,
  input  [1:0] io_cached_0_grant_bits_manager_xact_id,
  input   io_cached_0_grant_bits_is_builtin_type,
  input  [3:0] io_cached_0_grant_bits_g_type,
  input  [63:0] io_cached_0_grant_bits_data,
  input   io_cached_0_grant_bits_manager_id,
  input   io_cached_0_finish_ready,
  output  io_cached_0_finish_valid,
  output [1:0] io_cached_0_finish_bits_manager_xact_id,
  output  io_cached_0_finish_bits_manager_id,
  input   io_uncached_0_acquire_ready,
  output  io_uncached_0_acquire_valid,
  output [25:0] io_uncached_0_acquire_bits_addr_block,
  output  io_uncached_0_acquire_bits_client_xact_id,
  output [2:0] io_uncached_0_acquire_bits_addr_beat,
  output  io_uncached_0_acquire_bits_is_builtin_type,
  output [2:0] io_uncached_0_acquire_bits_a_type,
  output [11:0] io_uncached_0_acquire_bits_union,
  output [63:0] io_uncached_0_acquire_bits_data,
  output  io_uncached_0_grant_ready,
  input   io_uncached_0_grant_valid,
  input  [2:0] io_uncached_0_grant_bits_addr_beat,
  input   io_uncached_0_grant_bits_client_xact_id,
  input  [1:0] io_uncached_0_grant_bits_manager_xact_id,
  input   io_uncached_0_grant_bits_is_builtin_type,
  input  [3:0] io_uncached_0_grant_bits_g_type,
  input  [63:0] io_uncached_0_grant_bits_data,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip
);
//<CJ> RESET_VECTOR_ADDR
  parameter RESET_VECTOR_ADDR = 60000000;

  wire  core_clk;
  wire  core_reset;
  wire  core_io_prci_reset;
  wire  core_io_prci_id;
  wire  core_io_prci_interrupts_meip;
  wire  core_io_prci_interrupts_seip;
  wire  core_io_prci_interrupts_debug;
  wire  core_io_prci_interrupts_mtip;
  wire  core_io_prci_interrupts_msip;
  wire  core_io_imem_req_valid;
  wire [31:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_req_bits_speculative;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire [31:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data_0;
  wire  core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_if;
  wire  core_io_imem_resp_bits_replay;
  wire  core_io_imem_btb_resp_valid;
  wire  core_io_imem_btb_resp_bits_taken;
  wire  core_io_imem_btb_resp_bits_mask;
  wire  core_io_imem_btb_resp_bits_bridx;
  wire [31:0] core_io_imem_btb_resp_bits_target;
  wire  core_io_imem_btb_resp_bits_entry;
  wire  core_io_imem_btb_resp_bits_bht_history;
  wire [1:0] core_io_imem_btb_resp_bits_bht_value;
  wire  core_io_imem_btb_update_valid;
  wire  core_io_imem_btb_update_bits_prediction_valid;
  wire  core_io_imem_btb_update_bits_prediction_bits_taken;
  wire  core_io_imem_btb_update_bits_prediction_bits_mask;
  wire  core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire [31:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire  core_io_imem_btb_update_bits_prediction_bits_entry;
  wire  core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire [31:0] core_io_imem_btb_update_bits_pc;
  wire [31:0] core_io_imem_btb_update_bits_target;
  wire  core_io_imem_btb_update_bits_taken;
  wire  core_io_imem_btb_update_bits_isJump;
  wire  core_io_imem_btb_update_bits_isReturn;
  wire [31:0] core_io_imem_btb_update_bits_br_pc;
  wire  core_io_imem_bht_update_valid;
  wire  core_io_imem_bht_update_bits_prediction_valid;
  wire  core_io_imem_bht_update_bits_prediction_bits_taken;
  wire  core_io_imem_bht_update_bits_prediction_bits_mask;
  wire  core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire [31:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire  core_io_imem_bht_update_bits_prediction_bits_entry;
  wire  core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire [31:0] core_io_imem_bht_update_bits_pc;
  wire  core_io_imem_bht_update_bits_taken;
  wire  core_io_imem_bht_update_bits_mispredict;
  wire  core_io_imem_ras_update_valid;
  wire  core_io_imem_ras_update_bits_isCall;
  wire  core_io_imem_ras_update_bits_isReturn;
  wire [31:0] core_io_imem_ras_update_bits_returnAddr;
  wire  core_io_imem_ras_update_bits_prediction_valid;
  wire  core_io_imem_ras_update_bits_prediction_bits_taken;
  wire  core_io_imem_ras_update_bits_prediction_bits_mask;
  wire  core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire [31:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire  core_io_imem_ras_update_bits_prediction_bits_entry;
  wire  core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_flush_tlb;
  wire [31:0] core_io_imem_npc;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [31:0] core_io_dmem_req_bits_addr;
  wire [8:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire [31:0] core_io_dmem_req_bits_data;
  wire  core_io_dmem_s1_kill;
  wire [31:0] core_io_dmem_s1_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [31:0] core_io_dmem_resp_bits_addr;
  wire [8:0] core_io_dmem_resp_bits_tag;
  wire [4:0] core_io_dmem_resp_bits_cmd;
  wire [2:0] core_io_dmem_resp_bits_typ;
  wire [31:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [31:0] core_io_dmem_resp_bits_data_word_bypass;
  wire [31:0] core_io_dmem_resp_bits_store_data;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_xcpt_ma_ld;
  wire  core_io_dmem_xcpt_ma_st;
  wire  core_io_dmem_xcpt_pf_ld;
  wire  core_io_dmem_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [6:0] core_io_ptw_ptbr_asid;
  wire [21:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_invalidate;
  wire  core_io_ptw_status_debug;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_sd;
  wire [30:0] core_io_ptw_status_zero3;
  wire  core_io_ptw_status_sd_rv32;
  wire [1:0] core_io_ptw_status_zero2;
  wire [4:0] core_io_ptw_status_vm;
  wire [3:0] core_io_ptw_status_zero1;
  wire  core_io_ptw_status_mxr;
  wire  core_io_ptw_status_pum;
  wire  core_io_ptw_status_mprv;
  wire [1:0] core_io_ptw_status_xs;
  wire [1:0] core_io_ptw_status_fs;
  wire [1:0] core_io_ptw_status_mpp;
  wire [1:0] core_io_ptw_status_hpp;
  wire  core_io_ptw_status_spp;
  wire  core_io_ptw_status_mpie;
  wire  core_io_ptw_status_hpie;
  wire  core_io_ptw_status_spie;
  wire  core_io_ptw_status_upie;
  wire  core_io_ptw_status_mie;
  wire  core_io_ptw_status_hie;
  wire  core_io_ptw_status_sie;
  wire  core_io_ptw_status_uie;
  wire [31:0] core_io_fpu_inst;
  wire [31:0] core_io_fpu_fromint_data;
  wire [2:0] core_io_fpu_fcsr_rm;
  wire  core_io_fpu_fcsr_flags_valid;
  wire [4:0] core_io_fpu_fcsr_flags_bits;
  wire [63:0] core_io_fpu_store_data;
  wire [31:0] core_io_fpu_toint_data;
  wire  core_io_fpu_dmem_resp_val;
  wire [2:0] core_io_fpu_dmem_resp_type;
  wire [4:0] core_io_fpu_dmem_resp_tag;
  wire [63:0] core_io_fpu_dmem_resp_data;
  wire  core_io_fpu_valid;
  wire  core_io_fpu_fcsr_rdy;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_illegal_rm;
  wire  core_io_fpu_killx;
  wire  core_io_fpu_killm;
  wire [4:0] core_io_fpu_dec_cmd;
  wire  core_io_fpu_dec_ldst;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_fpu_dec_swap12;
  wire  core_io_fpu_dec_swap23;
  wire  core_io_fpu_dec_single;
  wire  core_io_fpu_dec_fromint;
  wire  core_io_fpu_dec_toint;
  wire  core_io_fpu_dec_fastpipe;
  wire  core_io_fpu_dec_fma;
  wire  core_io_fpu_dec_div;
  wire  core_io_fpu_dec_sqrt;
  wire  core_io_fpu_dec_round;
  wire  core_io_fpu_dec_wflags;
  wire  core_io_fpu_sboard_set;
  wire  core_io_fpu_sboard_clr;
  wire [4:0] core_io_fpu_sboard_clra;
  wire  core_io_fpu_cp_req_ready;
  wire  core_io_fpu_cp_req_valid;
  wire [4:0] core_io_fpu_cp_req_bits_cmd;
  wire  core_io_fpu_cp_req_bits_ldst;
  wire  core_io_fpu_cp_req_bits_wen;
  wire  core_io_fpu_cp_req_bits_ren1;
  wire  core_io_fpu_cp_req_bits_ren2;
  wire  core_io_fpu_cp_req_bits_ren3;
  wire  core_io_fpu_cp_req_bits_swap12;
  wire  core_io_fpu_cp_req_bits_swap23;
  wire  core_io_fpu_cp_req_bits_single;
  wire  core_io_fpu_cp_req_bits_fromint;
  wire  core_io_fpu_cp_req_bits_toint;
  wire  core_io_fpu_cp_req_bits_fastpipe;
  wire  core_io_fpu_cp_req_bits_fma;
  wire  core_io_fpu_cp_req_bits_div;
  wire  core_io_fpu_cp_req_bits_sqrt;
  wire  core_io_fpu_cp_req_bits_round;
  wire  core_io_fpu_cp_req_bits_wflags;
  wire [2:0] core_io_fpu_cp_req_bits_rm;
  wire [1:0] core_io_fpu_cp_req_bits_typ;
  wire [64:0] core_io_fpu_cp_req_bits_in1;
  wire [64:0] core_io_fpu_cp_req_bits_in2;
  wire [64:0] core_io_fpu_cp_req_bits_in3;
  wire  core_io_fpu_cp_resp_ready;
  wire  core_io_fpu_cp_resp_valid;
  wire [64:0] core_io_fpu_cp_resp_bits_data;
  wire [4:0] core_io_fpu_cp_resp_bits_exc;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_cmd_valid;
  wire [6:0] core_io_rocc_cmd_bits_inst_funct;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire  core_io_rocc_cmd_bits_inst_xd;
  wire  core_io_rocc_cmd_bits_inst_xs1;
  wire  core_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rd;
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire [31:0] core_io_rocc_cmd_bits_rs1;
  wire [31:0] core_io_rocc_cmd_bits_rs2;
  wire  core_io_rocc_cmd_bits_status_debug;
  wire [1:0] core_io_rocc_cmd_bits_status_prv;
  wire  core_io_rocc_cmd_bits_status_sd;
  wire [30:0] core_io_rocc_cmd_bits_status_zero3;
  wire  core_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] core_io_rocc_cmd_bits_status_zero2;
  wire [4:0] core_io_rocc_cmd_bits_status_vm;
  wire [3:0] core_io_rocc_cmd_bits_status_zero1;
  wire  core_io_rocc_cmd_bits_status_mxr;
  wire  core_io_rocc_cmd_bits_status_pum;
  wire  core_io_rocc_cmd_bits_status_mprv;
  wire [1:0] core_io_rocc_cmd_bits_status_xs;
  wire [1:0] core_io_rocc_cmd_bits_status_fs;
  wire [1:0] core_io_rocc_cmd_bits_status_mpp;
  wire [1:0] core_io_rocc_cmd_bits_status_hpp;
  wire  core_io_rocc_cmd_bits_status_spp;
  wire  core_io_rocc_cmd_bits_status_mpie;
  wire  core_io_rocc_cmd_bits_status_hpie;
  wire  core_io_rocc_cmd_bits_status_spie;
  wire  core_io_rocc_cmd_bits_status_upie;
  wire  core_io_rocc_cmd_bits_status_mie;
  wire  core_io_rocc_cmd_bits_status_hie;
  wire  core_io_rocc_cmd_bits_status_sie;
  wire  core_io_rocc_cmd_bits_status_uie;
  wire  core_io_rocc_resp_ready;
  wire  core_io_rocc_resp_valid;
  wire [4:0] core_io_rocc_resp_bits_rd;
  wire [31:0] core_io_rocc_resp_bits_data;
  wire  core_io_rocc_mem_req_ready;
  wire  core_io_rocc_mem_req_valid;
  wire [31:0] core_io_rocc_mem_req_bits_addr;
  wire [8:0] core_io_rocc_mem_req_bits_tag;
  wire [4:0] core_io_rocc_mem_req_bits_cmd;
  wire [2:0] core_io_rocc_mem_req_bits_typ;
  wire  core_io_rocc_mem_req_bits_phys;
  wire [31:0] core_io_rocc_mem_req_bits_data;
  wire  core_io_rocc_mem_s1_kill;
  wire [31:0] core_io_rocc_mem_s1_data;
  wire  core_io_rocc_mem_s2_nack;
  wire  core_io_rocc_mem_resp_valid;
  wire [31:0] core_io_rocc_mem_resp_bits_addr;
  wire [8:0] core_io_rocc_mem_resp_bits_tag;
  wire [4:0] core_io_rocc_mem_resp_bits_cmd;
  wire [2:0] core_io_rocc_mem_resp_bits_typ;
  wire [31:0] core_io_rocc_mem_resp_bits_data;
  wire  core_io_rocc_mem_resp_bits_replay;
  wire  core_io_rocc_mem_resp_bits_has_data;
  wire [31:0] core_io_rocc_mem_resp_bits_data_word_bypass;
  wire [31:0] core_io_rocc_mem_resp_bits_store_data;
  wire  core_io_rocc_mem_replay_next;
  wire  core_io_rocc_mem_xcpt_ma_ld;
  wire  core_io_rocc_mem_xcpt_ma_st;
  wire  core_io_rocc_mem_xcpt_pf_ld;
  wire  core_io_rocc_mem_xcpt_pf_st;
  wire  core_io_rocc_mem_invalidate_lr;
  wire  core_io_rocc_mem_ordered;
  wire  core_io_rocc_busy;
  wire  core_io_rocc_interrupt;
  wire  core_io_rocc_autl_acquire_ready;
  wire  core_io_rocc_autl_acquire_valid;
  wire [25:0] core_io_rocc_autl_acquire_bits_addr_block;
  wire  core_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_acquire_bits_addr_beat;
  wire  core_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] core_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] core_io_rocc_autl_acquire_bits_union;
  wire [63:0] core_io_rocc_autl_acquire_bits_data;
  wire  core_io_rocc_autl_grant_ready;
  wire  core_io_rocc_autl_grant_valid;
  wire [2:0] core_io_rocc_autl_grant_bits_addr_beat;
  wire  core_io_rocc_autl_grant_bits_client_xact_id;
  wire [1:0] core_io_rocc_autl_grant_bits_manager_xact_id;
  wire  core_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] core_io_rocc_autl_grant_bits_g_type;
  wire [63:0] core_io_rocc_autl_grant_bits_data;
  wire  core_io_rocc_fpu_req_ready;
  wire  core_io_rocc_fpu_req_valid;
  wire [4:0] core_io_rocc_fpu_req_bits_cmd;
  wire  core_io_rocc_fpu_req_bits_ldst;
  wire  core_io_rocc_fpu_req_bits_wen;
  wire  core_io_rocc_fpu_req_bits_ren1;
  wire  core_io_rocc_fpu_req_bits_ren2;
  wire  core_io_rocc_fpu_req_bits_ren3;
  wire  core_io_rocc_fpu_req_bits_swap12;
  wire  core_io_rocc_fpu_req_bits_swap23;
  wire  core_io_rocc_fpu_req_bits_single;
  wire  core_io_rocc_fpu_req_bits_fromint;
  wire  core_io_rocc_fpu_req_bits_toint;
  wire  core_io_rocc_fpu_req_bits_fastpipe;
  wire  core_io_rocc_fpu_req_bits_fma;
  wire  core_io_rocc_fpu_req_bits_div;
  wire  core_io_rocc_fpu_req_bits_sqrt;
  wire  core_io_rocc_fpu_req_bits_round;
  wire  core_io_rocc_fpu_req_bits_wflags;
  wire [2:0] core_io_rocc_fpu_req_bits_rm;
  wire [1:0] core_io_rocc_fpu_req_bits_typ;
  wire [64:0] core_io_rocc_fpu_req_bits_in1;
  wire [64:0] core_io_rocc_fpu_req_bits_in2;
  wire [64:0] core_io_rocc_fpu_req_bits_in3;
  wire  core_io_rocc_fpu_resp_ready;
  wire  core_io_rocc_fpu_resp_valid;
  wire [64:0] core_io_rocc_fpu_resp_bits_data;
  wire [4:0] core_io_rocc_fpu_resp_bits_exc;
  wire  core_io_rocc_exception;
  wire [11:0] core_io_rocc_csr_waddr;
  wire [31:0] core_io_rocc_csr_wdata;
  wire  core_io_rocc_csr_wen;
  wire  core_io_rocc_host_id;
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_cpu_req_valid;
  wire [31:0] icache_io_cpu_req_bits_pc;
  wire  icache_io_cpu_req_bits_speculative;
  wire  icache_io_cpu_resp_ready;
  wire  icache_io_cpu_resp_valid;
  wire [31:0] icache_io_cpu_resp_bits_pc;
  wire [31:0] icache_io_cpu_resp_bits_data_0;
  wire  icache_io_cpu_resp_bits_mask;
  wire  icache_io_cpu_resp_bits_xcpt_if;
  wire  icache_io_cpu_resp_bits_replay;
  wire  icache_io_cpu_btb_resp_valid;
  wire  icache_io_cpu_btb_resp_bits_taken;
  wire  icache_io_cpu_btb_resp_bits_mask;
  wire  icache_io_cpu_btb_resp_bits_bridx;
  wire [31:0] icache_io_cpu_btb_resp_bits_target;
  wire  icache_io_cpu_btb_resp_bits_entry;
  wire  icache_io_cpu_btb_resp_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire  icache_io_cpu_btb_update_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bridx;
  wire [31:0] icache_io_cpu_btb_update_bits_prediction_bits_target;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_value;
  wire [31:0] icache_io_cpu_btb_update_bits_pc;
  wire [31:0] icache_io_cpu_btb_update_bits_target;
  wire  icache_io_cpu_btb_update_bits_taken;
  wire  icache_io_cpu_btb_update_bits_isJump;
  wire  icache_io_cpu_btb_update_bits_isReturn;
  wire [31:0] icache_io_cpu_btb_update_bits_br_pc;
  wire  icache_io_cpu_bht_update_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bridx;
  wire [31:0] icache_io_cpu_bht_update_bits_prediction_bits_target;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_value;
  wire [31:0] icache_io_cpu_bht_update_bits_pc;
  wire  icache_io_cpu_bht_update_bits_taken;
  wire  icache_io_cpu_bht_update_bits_mispredict;
  wire  icache_io_cpu_ras_update_valid;
  wire  icache_io_cpu_ras_update_bits_isCall;
  wire  icache_io_cpu_ras_update_bits_isReturn;
  wire [31:0] icache_io_cpu_ras_update_bits_returnAddr;
  wire  icache_io_cpu_ras_update_bits_prediction_valid;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bridx;
  wire [31:0] icache_io_cpu_ras_update_bits_prediction_bits_target;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_value;
  wire  icache_io_cpu_flush_icache;
  wire  icache_io_cpu_flush_tlb;
  wire [31:0] icache_io_cpu_npc;
  wire  icache_io_ptw_req_ready;
  wire  icache_io_ptw_req_valid;
  wire [1:0] icache_io_ptw_req_bits_prv;
  wire  icache_io_ptw_req_bits_pum;
  wire  icache_io_ptw_req_bits_mxr;
  wire [19:0] icache_io_ptw_req_bits_addr;
  wire  icache_io_ptw_req_bits_store;
  wire  icache_io_ptw_req_bits_fetch;
  wire  icache_io_ptw_resp_valid;
  wire [15:0] icache_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] icache_io_ptw_resp_bits_pte_ppn;
  wire [1:0] icache_io_ptw_resp_bits_pte_reserved_for_software;
  wire  icache_io_ptw_resp_bits_pte_d;
  wire  icache_io_ptw_resp_bits_pte_a;
  wire  icache_io_ptw_resp_bits_pte_g;
  wire  icache_io_ptw_resp_bits_pte_u;
  wire  icache_io_ptw_resp_bits_pte_x;
  wire  icache_io_ptw_resp_bits_pte_w;
  wire  icache_io_ptw_resp_bits_pte_r;
  wire  icache_io_ptw_resp_bits_pte_v;
  wire [6:0] icache_io_ptw_ptbr_asid;
  wire [21:0] icache_io_ptw_ptbr_ppn;
  wire  icache_io_ptw_invalidate;
  wire  icache_io_ptw_status_debug;
  wire [1:0] icache_io_ptw_status_prv;
  wire  icache_io_ptw_status_sd;
  wire [30:0] icache_io_ptw_status_zero3;
  wire  icache_io_ptw_status_sd_rv32;
  wire [1:0] icache_io_ptw_status_zero2;
  wire [4:0] icache_io_ptw_status_vm;
  wire [3:0] icache_io_ptw_status_zero1;
  wire  icache_io_ptw_status_mxr;
  wire  icache_io_ptw_status_pum;
  wire  icache_io_ptw_status_mprv;
  wire [1:0] icache_io_ptw_status_xs;
  wire [1:0] icache_io_ptw_status_fs;
  wire [1:0] icache_io_ptw_status_mpp;
  wire [1:0] icache_io_ptw_status_hpp;
  wire  icache_io_ptw_status_spp;
  wire  icache_io_ptw_status_mpie;
  wire  icache_io_ptw_status_hpie;
  wire  icache_io_ptw_status_spie;
  wire  icache_io_ptw_status_upie;
  wire  icache_io_ptw_status_mie;
  wire  icache_io_ptw_status_hie;
  wire  icache_io_ptw_status_sie;
  wire  icache_io_ptw_status_uie;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire  icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire  icache_io_mem_grant_bits_client_xact_id;
  wire [1:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  DCache_1_clk;
  wire  DCache_1_reset;
  wire  DCache_1_io_cpu_req_ready;
  wire  DCache_1_io_cpu_req_valid;
  wire [31:0] DCache_1_io_cpu_req_bits_addr;
  wire [8:0] DCache_1_io_cpu_req_bits_tag;
  wire [4:0] DCache_1_io_cpu_req_bits_cmd;
  wire [2:0] DCache_1_io_cpu_req_bits_typ;
  wire  DCache_1_io_cpu_req_bits_phys;
  wire [31:0] DCache_1_io_cpu_req_bits_data;
  wire  DCache_1_io_cpu_s1_kill;
  wire [31:0] DCache_1_io_cpu_s1_data;
  wire  DCache_1_io_cpu_s2_nack;
  wire  DCache_1_io_cpu_resp_valid;
  wire [31:0] DCache_1_io_cpu_resp_bits_addr;
  wire [8:0] DCache_1_io_cpu_resp_bits_tag;
  wire [4:0] DCache_1_io_cpu_resp_bits_cmd;
  wire [2:0] DCache_1_io_cpu_resp_bits_typ;
  wire [31:0] DCache_1_io_cpu_resp_bits_data;
  wire  DCache_1_io_cpu_resp_bits_replay;
  wire  DCache_1_io_cpu_resp_bits_has_data;
  wire [31:0] DCache_1_io_cpu_resp_bits_data_word_bypass;
  wire [31:0] DCache_1_io_cpu_resp_bits_store_data;
  wire  DCache_1_io_cpu_replay_next;
  wire  DCache_1_io_cpu_xcpt_ma_ld;
  wire  DCache_1_io_cpu_xcpt_ma_st;
  wire  DCache_1_io_cpu_xcpt_pf_ld;
  wire  DCache_1_io_cpu_xcpt_pf_st;
  wire  DCache_1_io_cpu_invalidate_lr;
  wire  DCache_1_io_cpu_ordered;
  wire  DCache_1_io_ptw_req_ready;
  wire  DCache_1_io_ptw_req_valid;
  wire [1:0] DCache_1_io_ptw_req_bits_prv;
  wire  DCache_1_io_ptw_req_bits_pum;
  wire  DCache_1_io_ptw_req_bits_mxr;
  wire [19:0] DCache_1_io_ptw_req_bits_addr;
  wire  DCache_1_io_ptw_req_bits_store;
  wire  DCache_1_io_ptw_req_bits_fetch;
  wire  DCache_1_io_ptw_resp_valid;
  wire [15:0] DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] DCache_1_io_ptw_resp_bits_pte_ppn;
  wire [1:0] DCache_1_io_ptw_resp_bits_pte_reserved_for_software;
  wire  DCache_1_io_ptw_resp_bits_pte_d;
  wire  DCache_1_io_ptw_resp_bits_pte_a;
  wire  DCache_1_io_ptw_resp_bits_pte_g;
  wire  DCache_1_io_ptw_resp_bits_pte_u;
  wire  DCache_1_io_ptw_resp_bits_pte_x;
  wire  DCache_1_io_ptw_resp_bits_pte_w;
  wire  DCache_1_io_ptw_resp_bits_pte_r;
  wire  DCache_1_io_ptw_resp_bits_pte_v;
  wire [6:0] DCache_1_io_ptw_ptbr_asid;
  wire [21:0] DCache_1_io_ptw_ptbr_ppn;
  wire  DCache_1_io_ptw_invalidate;
  wire  DCache_1_io_ptw_status_debug;
  wire [1:0] DCache_1_io_ptw_status_prv;
  wire  DCache_1_io_ptw_status_sd;
  wire [30:0] DCache_1_io_ptw_status_zero3;
  wire  DCache_1_io_ptw_status_sd_rv32;
  wire [1:0] DCache_1_io_ptw_status_zero2;
  wire [4:0] DCache_1_io_ptw_status_vm;
  wire [3:0] DCache_1_io_ptw_status_zero1;
  wire  DCache_1_io_ptw_status_mxr;
  wire  DCache_1_io_ptw_status_pum;
  wire  DCache_1_io_ptw_status_mprv;
  wire [1:0] DCache_1_io_ptw_status_xs;
  wire [1:0] DCache_1_io_ptw_status_fs;
  wire [1:0] DCache_1_io_ptw_status_mpp;
  wire [1:0] DCache_1_io_ptw_status_hpp;
  wire  DCache_1_io_ptw_status_spp;
  wire  DCache_1_io_ptw_status_mpie;
  wire  DCache_1_io_ptw_status_hpie;
  wire  DCache_1_io_ptw_status_spie;
  wire  DCache_1_io_ptw_status_upie;
  wire  DCache_1_io_ptw_status_mie;
  wire  DCache_1_io_ptw_status_hie;
  wire  DCache_1_io_ptw_status_sie;
  wire  DCache_1_io_ptw_status_uie;
  wire  DCache_1_io_mem_acquire_ready;
  wire  DCache_1_io_mem_acquire_valid;
  wire [25:0] DCache_1_io_mem_acquire_bits_addr_block;
  wire  DCache_1_io_mem_acquire_bits_client_xact_id;
  wire [2:0] DCache_1_io_mem_acquire_bits_addr_beat;
  wire  DCache_1_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] DCache_1_io_mem_acquire_bits_a_type;
  wire [11:0] DCache_1_io_mem_acquire_bits_union;
  wire [63:0] DCache_1_io_mem_acquire_bits_data;
  wire  DCache_1_io_mem_probe_ready;
  wire  DCache_1_io_mem_probe_valid;
  wire [25:0] DCache_1_io_mem_probe_bits_addr_block;
  wire [1:0] DCache_1_io_mem_probe_bits_p_type;
  wire  DCache_1_io_mem_release_ready;
  wire  DCache_1_io_mem_release_valid;
  wire [2:0] DCache_1_io_mem_release_bits_addr_beat;
  wire [25:0] DCache_1_io_mem_release_bits_addr_block;
  wire  DCache_1_io_mem_release_bits_client_xact_id;
  wire  DCache_1_io_mem_release_bits_voluntary;
  wire [2:0] DCache_1_io_mem_release_bits_r_type;
  wire [63:0] DCache_1_io_mem_release_bits_data;
  wire  DCache_1_io_mem_grant_ready;
  wire  DCache_1_io_mem_grant_valid;
  wire [2:0] DCache_1_io_mem_grant_bits_addr_beat;
  wire  DCache_1_io_mem_grant_bits_client_xact_id;
  wire [1:0] DCache_1_io_mem_grant_bits_manager_xact_id;
  wire  DCache_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] DCache_1_io_mem_grant_bits_g_type;
  wire [63:0] DCache_1_io_mem_grant_bits_data;
  wire  DCache_1_io_mem_grant_bits_manager_id;
  wire  DCache_1_io_mem_finish_ready;
  wire  DCache_1_io_mem_finish_valid;
  wire [1:0] DCache_1_io_mem_finish_bits_manager_xact_id;
  wire  DCache_1_io_mem_finish_bits_manager_id;
  wire  uncachedArb_clk;
  wire  uncachedArb_reset;
  wire  uncachedArb_io_in_0_acquire_ready;
  wire  uncachedArb_io_in_0_acquire_valid;
  wire [25:0] uncachedArb_io_in_0_acquire_bits_addr_block;
  wire  uncachedArb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_addr_beat;
  wire  uncachedArb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_in_0_acquire_bits_union;
  wire [63:0] uncachedArb_io_in_0_acquire_bits_data;
  wire  uncachedArb_io_in_0_grant_ready;
  wire  uncachedArb_io_in_0_grant_valid;
  wire [2:0] uncachedArb_io_in_0_grant_bits_addr_beat;
  wire  uncachedArb_io_in_0_grant_bits_client_xact_id;
  wire [1:0] uncachedArb_io_in_0_grant_bits_manager_xact_id;
  wire  uncachedArb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_in_0_grant_bits_g_type;
  wire [63:0] uncachedArb_io_in_0_grant_bits_data;
  wire  uncachedArb_io_out_acquire_ready;
  wire  uncachedArb_io_out_acquire_valid;
  wire [25:0] uncachedArb_io_out_acquire_bits_addr_block;
  wire  uncachedArb_io_out_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_acquire_bits_addr_beat;
  wire  uncachedArb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_out_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_out_acquire_bits_union;
  wire [63:0] uncachedArb_io_out_acquire_bits_data;
  wire  uncachedArb_io_out_grant_ready;
  wire  uncachedArb_io_out_grant_valid;
  wire [2:0] uncachedArb_io_out_grant_bits_addr_beat;
  wire  uncachedArb_io_out_grant_bits_client_xact_id;
  wire [1:0] uncachedArb_io_out_grant_bits_manager_xact_id;
  wire  uncachedArb_io_out_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_out_grant_bits_g_type;
  wire [63:0] uncachedArb_io_out_grant_bits_data;
  wire  dcArb_clk;
  wire  dcArb_reset;
  wire  dcArb_io_requestor_0_req_ready;
  wire  dcArb_io_requestor_0_req_valid;
  wire [31:0] dcArb_io_requestor_0_req_bits_addr;
  wire [8:0] dcArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_req_bits_typ;
  wire  dcArb_io_requestor_0_req_bits_phys;
  wire [31:0] dcArb_io_requestor_0_req_bits_data;
  wire  dcArb_io_requestor_0_s1_kill;
  wire [31:0] dcArb_io_requestor_0_s1_data;
  wire  dcArb_io_requestor_0_s2_nack;
  wire  dcArb_io_requestor_0_resp_valid;
  wire [31:0] dcArb_io_requestor_0_resp_bits_addr;
  wire [8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire [31:0] dcArb_io_requestor_0_resp_bits_data;
  wire  dcArb_io_requestor_0_resp_bits_replay;
  wire  dcArb_io_requestor_0_resp_bits_has_data;
  wire [31:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire [31:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire  dcArb_io_requestor_0_replay_next;
  wire  dcArb_io_requestor_0_xcpt_ma_ld;
  wire  dcArb_io_requestor_0_xcpt_ma_st;
  wire  dcArb_io_requestor_0_xcpt_pf_ld;
  wire  dcArb_io_requestor_0_xcpt_pf_st;
  wire  dcArb_io_requestor_0_invalidate_lr;
  wire  dcArb_io_requestor_0_ordered;
  wire  dcArb_io_mem_req_ready;
  wire  dcArb_io_mem_req_valid;
  wire [31:0] dcArb_io_mem_req_bits_addr;
  wire [8:0] dcArb_io_mem_req_bits_tag;
  wire [4:0] dcArb_io_mem_req_bits_cmd;
  wire [2:0] dcArb_io_mem_req_bits_typ;
  wire  dcArb_io_mem_req_bits_phys;
  wire [31:0] dcArb_io_mem_req_bits_data;
  wire  dcArb_io_mem_s1_kill;
  wire [31:0] dcArb_io_mem_s1_data;
  wire  dcArb_io_mem_s2_nack;
  wire  dcArb_io_mem_resp_valid;
  wire [31:0] dcArb_io_mem_resp_bits_addr;
  wire [8:0] dcArb_io_mem_resp_bits_tag;
  wire [4:0] dcArb_io_mem_resp_bits_cmd;
  wire [2:0] dcArb_io_mem_resp_bits_typ;
  wire [31:0] dcArb_io_mem_resp_bits_data;
  wire  dcArb_io_mem_resp_bits_replay;
  wire  dcArb_io_mem_resp_bits_has_data;
  wire [31:0] dcArb_io_mem_resp_bits_data_word_bypass;
  wire [31:0] dcArb_io_mem_resp_bits_store_data;
  wire  dcArb_io_mem_replay_next;
  wire  dcArb_io_mem_xcpt_ma_ld;
  wire  dcArb_io_mem_xcpt_ma_st;
  wire  dcArb_io_mem_xcpt_pf_ld;
  wire  dcArb_io_mem_xcpt_pf_st;
  wire  dcArb_io_mem_invalidate_lr;
  wire  dcArb_io_mem_ordered;
  reg  GEN_0;
  reg [31:0] GEN_160;
  reg [4:0] GEN_1;
  reg [31:0] GEN_161;
  reg [63:0] GEN_2;
  reg [63:0] GEN_162;
  reg [31:0] GEN_3;
  reg [31:0] GEN_163;
  reg  GEN_4;
  reg [31:0] GEN_164;
  reg  GEN_5;
  reg [31:0] GEN_165;
  reg  GEN_6;
  reg [31:0] GEN_166;
  reg [4:0] GEN_7;
  reg [31:0] GEN_167;
  reg  GEN_8;
  reg [31:0] GEN_168;
  reg  GEN_9;
  reg [31:0] GEN_169;
  reg  GEN_10;
  reg [31:0] GEN_170;
  reg  GEN_11;
  reg [31:0] GEN_171;
  reg  GEN_12;
  reg [31:0] GEN_172;
  reg  GEN_13;
  reg [31:0] GEN_173;
  reg  GEN_14;
  reg [31:0] GEN_174;
  reg  GEN_15;
  reg [31:0] GEN_175;
  reg  GEN_16;
  reg [31:0] GEN_176;
  reg  GEN_17;
  reg [31:0] GEN_177;
  reg  GEN_18;
  reg [31:0] GEN_178;
  reg  GEN_19;
  reg [31:0] GEN_179;
  reg  GEN_20;
  reg [31:0] GEN_180;
  reg  GEN_21;
  reg [31:0] GEN_181;
  reg  GEN_22;
  reg [31:0] GEN_182;
  reg  GEN_23;
  reg [31:0] GEN_183;
  reg  GEN_24;
  reg [31:0] GEN_184;
  reg  GEN_25;
  reg [31:0] GEN_185;
  reg [4:0] GEN_26;
  reg [31:0] GEN_186;
  reg  GEN_27;
  reg [31:0] GEN_187;
  reg  GEN_28;
  reg [31:0] GEN_188;
  reg [64:0] GEN_29;
  reg [95:0] GEN_189;
  reg [4:0] GEN_30;
  reg [31:0] GEN_190;
  reg  GEN_31;
  reg [31:0] GEN_191;
  reg  GEN_32;
  reg [31:0] GEN_192;
  reg [4:0] GEN_33;
  reg [31:0] GEN_193;
  reg [31:0] GEN_34;
  reg [31:0] GEN_194;
  reg  GEN_35;
  reg [31:0] GEN_195;
  reg [31:0] GEN_36;
  reg [31:0] GEN_196;
  reg [8:0] GEN_37;
  reg [31:0] GEN_197;
  reg [4:0] GEN_38;
  reg [31:0] GEN_198;
  reg [2:0] GEN_39;
  reg [31:0] GEN_199;
  reg  GEN_40;
  reg [31:0] GEN_200;
  reg [31:0] GEN_41;
  reg [31:0] GEN_201;
  reg  GEN_42;
  reg [31:0] GEN_202;
  reg [31:0] GEN_43;
  reg [31:0] GEN_203;
  reg  GEN_44;
  reg [31:0] GEN_204;
  reg  GEN_45;
  reg [31:0] GEN_205;
  reg  GEN_46;
  reg [31:0] GEN_206;
  reg  GEN_47;
  reg [31:0] GEN_207;
  reg [25:0] GEN_48;
  reg [31:0] GEN_208;
  reg  GEN_49;
  reg [31:0] GEN_209;
  reg [2:0] GEN_50;
  reg [31:0] GEN_210;
  reg  GEN_51;
  reg [31:0] GEN_211;
  reg [2:0] GEN_52;
  reg [31:0] GEN_212;
  reg [11:0] GEN_53;
  reg [31:0] GEN_213;
  reg [63:0] GEN_54;
  reg [63:0] GEN_214;
  reg  GEN_55;
  reg [31:0] GEN_215;
  reg  GEN_56;
  reg [31:0] GEN_216;
  reg [4:0] GEN_57;
  reg [31:0] GEN_217;
  reg  GEN_58;
  reg [31:0] GEN_218;
  reg  GEN_59;
  reg [31:0] GEN_219;
  reg  GEN_60;
  reg [31:0] GEN_220;
  reg  GEN_61;
  reg [31:0] GEN_221;
  reg  GEN_62;
  reg [31:0] GEN_222;
  reg  GEN_63;
  reg [31:0] GEN_223;
  reg  GEN_64;
  reg [31:0] GEN_224;
  reg  GEN_65;
  reg [31:0] GEN_225;
  reg  GEN_66;
  reg [31:0] GEN_226;
  reg  GEN_67;
  reg [31:0] GEN_227;
  reg  GEN_68;
  reg [31:0] GEN_228;
  reg  GEN_69;
  reg [31:0] GEN_229;
  reg  GEN_70;
  reg [31:0] GEN_230;
  reg  GEN_71;
  reg [31:0] GEN_231;
  reg  GEN_72;
  reg [31:0] GEN_232;
  reg  GEN_73;
  reg [31:0] GEN_233;
  reg [2:0] GEN_74;
  reg [31:0] GEN_234;
  reg [1:0] GEN_75;
  reg [31:0] GEN_235;
  reg [64:0] GEN_76;
  reg [95:0] GEN_236;
  reg [64:0] GEN_77;
  reg [95:0] GEN_237;
  reg [64:0] GEN_78;
  reg [95:0] GEN_238;
  reg  GEN_79;
  reg [31:0] GEN_239;
  reg  GEN_80;
  reg [31:0] GEN_240;
  reg  GEN_81;
  reg [31:0] GEN_241;
  reg [15:0] GEN_82;
  reg [31:0] GEN_242;
  reg [37:0] GEN_83;
  reg [63:0] GEN_243;
  reg [1:0] GEN_84;
  reg [31:0] GEN_244;
  reg  GEN_85;
  reg [31:0] GEN_245;
  reg  GEN_86;
  reg [31:0] GEN_246;
  reg  GEN_87;
  reg [31:0] GEN_247;
  reg  GEN_88;
  reg [31:0] GEN_248;
  reg  GEN_89;
  reg [31:0] GEN_249;
  reg  GEN_90;
  reg [31:0] GEN_250;
  reg  GEN_91;
  reg [31:0] GEN_251;
  reg  GEN_92;
  reg [31:0] GEN_252;
  reg [6:0] GEN_93;
  reg [31:0] GEN_253;
  reg [21:0] GEN_94;
  reg [31:0] GEN_254;
  reg  GEN_95;
  reg [31:0] GEN_255;
  reg  GEN_96;
  reg [31:0] GEN_256;
  reg [1:0] GEN_97;
  reg [31:0] GEN_257;
  reg  GEN_98;
  reg [31:0] GEN_258;
  reg [30:0] GEN_99;
  reg [31:0] GEN_259;
  reg  GEN_100;
  reg [31:0] GEN_260;
  reg [1:0] GEN_101;
  reg [31:0] GEN_261;
  reg [4:0] GEN_102;
  reg [31:0] GEN_262;
  reg [3:0] GEN_103;
  reg [31:0] GEN_263;
  reg  GEN_104;
  reg [31:0] GEN_264;
  reg  GEN_105;
  reg [31:0] GEN_265;
  reg  GEN_106;
  reg [31:0] GEN_266;
  reg [1:0] GEN_107;
  reg [31:0] GEN_267;
  reg [1:0] GEN_108;
  reg [31:0] GEN_268;
  reg [1:0] GEN_109;
  reg [31:0] GEN_269;
  reg [1:0] GEN_110;
  reg [31:0] GEN_270;
  reg  GEN_111;
  reg [31:0] GEN_271;
  reg  GEN_112;
  reg [31:0] GEN_272;
  reg  GEN_113;
  reg [31:0] GEN_273;
  reg  GEN_114;
  reg [31:0] GEN_274;
  reg  GEN_115;
  reg [31:0] GEN_275;
  reg  GEN_116;
  reg [31:0] GEN_276;
  reg  GEN_117;
  reg [31:0] GEN_277;
  reg  GEN_118;
  reg [31:0] GEN_278;
  reg  GEN_119;
  reg [31:0] GEN_279;
  reg  GEN_120;
  reg [31:0] GEN_280;
  reg  GEN_121;
  reg [31:0] GEN_281;
  reg [15:0] GEN_122;
  reg [31:0] GEN_282;
  reg [37:0] GEN_123;
  reg [63:0] GEN_283;
  reg [1:0] GEN_124;
  reg [31:0] GEN_284;
  reg  GEN_125;
  reg [31:0] GEN_285;
  reg  GEN_126;
  reg [31:0] GEN_286;
  reg  GEN_127;
  reg [31:0] GEN_287;
  reg  GEN_128;
  reg [31:0] GEN_288;
  reg  GEN_129;
  reg [31:0] GEN_289;
  reg  GEN_130;
  reg [31:0] GEN_290;
  reg  GEN_131;
  reg [31:0] GEN_291;
  reg  GEN_132;
  reg [31:0] GEN_292;
  reg [6:0] GEN_133;
  reg [31:0] GEN_293;
  reg [21:0] GEN_134;
  reg [31:0] GEN_294;
  reg  GEN_135;
  reg [31:0] GEN_295;
  reg  GEN_136;
  reg [31:0] GEN_296;
  reg [1:0] GEN_137;
  reg [31:0] GEN_297;
  reg  GEN_138;
  reg [31:0] GEN_298;
  reg [30:0] GEN_139;
  reg [31:0] GEN_299;
  reg  GEN_140;
  reg [31:0] GEN_300;
  reg [1:0] GEN_141;
  reg [31:0] GEN_301;
  reg [4:0] GEN_142;
  reg [31:0] GEN_302;
  reg [3:0] GEN_143;
  reg [31:0] GEN_303;
  reg  GEN_144;
  reg [31:0] GEN_304;
  reg  GEN_145;
  reg [31:0] GEN_305;
  reg  GEN_146;
  reg [31:0] GEN_306;
  reg [1:0] GEN_147;
  reg [31:0] GEN_307;
  reg [1:0] GEN_148;
  reg [31:0] GEN_308;
  reg [1:0] GEN_149;
  reg [31:0] GEN_309;
  reg [1:0] GEN_150;
  reg [31:0] GEN_310;
  reg  GEN_151;
  reg [31:0] GEN_311;
  reg  GEN_152;
  reg [31:0] GEN_312;
  reg  GEN_153;
  reg [31:0] GEN_313;
  reg  GEN_154;
  reg [31:0] GEN_314;
  reg  GEN_155;
  reg [31:0] GEN_315;
  reg  GEN_156;
  reg [31:0] GEN_316;
  reg  GEN_157;
  reg [31:0] GEN_317;
  reg  GEN_158;
  reg [31:0] GEN_318;
  reg  GEN_159;
  reg [31:0] GEN_319;
  CORERISCV_AXI4_ROCKET core (
    .clk(core_clk),
    .reset(core_reset),
    .io_prci_reset(core_io_prci_reset),
    .io_prci_id(core_io_prci_id),
    .io_prci_interrupts_meip(core_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(core_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(core_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(core_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(core_io_prci_interrupts_msip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data_0(core_io_imem_resp_bits_data_0),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_if(core_io_imem_resp_bits_xcpt_if),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_resp_valid(core_io_imem_btb_resp_valid),
    .io_imem_btb_resp_bits_taken(core_io_imem_btb_resp_bits_taken),
    .io_imem_btb_resp_bits_mask(core_io_imem_btb_resp_bits_mask),
    .io_imem_btb_resp_bits_bridx(core_io_imem_btb_resp_bits_bridx),
    .io_imem_btb_resp_bits_target(core_io_imem_btb_resp_bits_target),
    .io_imem_btb_resp_bits_entry(core_io_imem_btb_resp_bits_entry),
    .io_imem_btb_resp_bits_bht_history(core_io_imem_btb_resp_bits_bht_history),
    .io_imem_btb_resp_bits_bht_value(core_io_imem_btb_resp_bits_bht_value),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_valid(core_io_imem_btb_update_bits_prediction_valid),
    .io_imem_btb_update_bits_prediction_bits_taken(core_io_imem_btb_update_bits_prediction_bits_taken),
    .io_imem_btb_update_bits_prediction_bits_mask(core_io_imem_btb_update_bits_prediction_bits_mask),
    .io_imem_btb_update_bits_prediction_bits_bridx(core_io_imem_btb_update_bits_prediction_bits_bridx),
    .io_imem_btb_update_bits_prediction_bits_target(core_io_imem_btb_update_bits_prediction_bits_target),
    .io_imem_btb_update_bits_prediction_bits_entry(core_io_imem_btb_update_bits_prediction_bits_entry),
    .io_imem_btb_update_bits_prediction_bits_bht_history(core_io_imem_btb_update_bits_prediction_bits_bht_history),
    .io_imem_btb_update_bits_prediction_bits_bht_value(core_io_imem_btb_update_bits_prediction_bits_bht_value),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_target(core_io_imem_btb_update_bits_target),
    .io_imem_btb_update_bits_taken(core_io_imem_btb_update_bits_taken),
    .io_imem_btb_update_bits_isJump(core_io_imem_btb_update_bits_isJump),
    .io_imem_btb_update_bits_isReturn(core_io_imem_btb_update_bits_isReturn),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_valid(core_io_imem_bht_update_bits_prediction_valid),
    .io_imem_bht_update_bits_prediction_bits_taken(core_io_imem_bht_update_bits_prediction_bits_taken),
    .io_imem_bht_update_bits_prediction_bits_mask(core_io_imem_bht_update_bits_prediction_bits_mask),
    .io_imem_bht_update_bits_prediction_bits_bridx(core_io_imem_bht_update_bits_prediction_bits_bridx),
    .io_imem_bht_update_bits_prediction_bits_target(core_io_imem_bht_update_bits_prediction_bits_target),
    .io_imem_bht_update_bits_prediction_bits_entry(core_io_imem_bht_update_bits_prediction_bits_entry),
    .io_imem_bht_update_bits_prediction_bits_bht_history(core_io_imem_bht_update_bits_prediction_bits_bht_history),
    .io_imem_bht_update_bits_prediction_bits_bht_value(core_io_imem_bht_update_bits_prediction_bits_bht_value),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_ras_update_valid(core_io_imem_ras_update_valid),
    .io_imem_ras_update_bits_isCall(core_io_imem_ras_update_bits_isCall),
    .io_imem_ras_update_bits_isReturn(core_io_imem_ras_update_bits_isReturn),
    .io_imem_ras_update_bits_returnAddr(core_io_imem_ras_update_bits_returnAddr),
    .io_imem_ras_update_bits_prediction_valid(core_io_imem_ras_update_bits_prediction_valid),
    .io_imem_ras_update_bits_prediction_bits_taken(core_io_imem_ras_update_bits_prediction_bits_taken),
    .io_imem_ras_update_bits_prediction_bits_mask(core_io_imem_ras_update_bits_prediction_bits_mask),
    .io_imem_ras_update_bits_prediction_bits_bridx(core_io_imem_ras_update_bits_prediction_bits_bridx),
    .io_imem_ras_update_bits_prediction_bits_target(core_io_imem_ras_update_bits_prediction_bits_target),
    .io_imem_ras_update_bits_prediction_bits_entry(core_io_imem_ras_update_bits_prediction_bits_entry),
    .io_imem_ras_update_bits_prediction_bits_bht_history(core_io_imem_ras_update_bits_prediction_bits_bht_history),
    .io_imem_ras_update_bits_prediction_bits_bht_value(core_io_imem_ras_update_bits_prediction_bits_bht_value),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_flush_tlb(core_io_imem_flush_tlb),
    .io_imem_npc(core_io_imem_npc),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data(core_io_dmem_s1_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_addr(core_io_dmem_resp_bits_addr),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_cmd(core_io_dmem_resp_bits_cmd),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_resp_bits_store_data(core_io_dmem_resp_bits_store_data),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_xcpt_ma_ld(core_io_dmem_xcpt_ma_ld),
    .io_dmem_xcpt_ma_st(core_io_dmem_xcpt_ma_st),
    .io_dmem_xcpt_pf_ld(core_io_dmem_xcpt_pf_ld),
    .io_dmem_xcpt_pf_st(core_io_dmem_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr_asid(core_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(core_io_ptw_invalidate),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero3(core_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_vm(core_io_ptw_status_vm),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_pum(core_io_ptw_status_pum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_hpp(core_io_ptw_status_hpp),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_cmd(core_io_fpu_dec_cmd),
    .io_fpu_dec_ldst(core_io_fpu_dec_ldst),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_dec_swap12(core_io_fpu_dec_swap12),
    .io_fpu_dec_swap23(core_io_fpu_dec_swap23),
    .io_fpu_dec_single(core_io_fpu_dec_single),
    .io_fpu_dec_fromint(core_io_fpu_dec_fromint),
    .io_fpu_dec_toint(core_io_fpu_dec_toint),
    .io_fpu_dec_fastpipe(core_io_fpu_dec_fastpipe),
    .io_fpu_dec_fma(core_io_fpu_dec_fma),
    .io_fpu_dec_div(core_io_fpu_dec_div),
    .io_fpu_dec_sqrt(core_io_fpu_dec_sqrt),
    .io_fpu_dec_round(core_io_fpu_dec_round),
    .io_fpu_dec_wflags(core_io_fpu_dec_wflags),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_fpu_cp_req_ready(core_io_fpu_cp_req_ready),
    .io_fpu_cp_req_valid(core_io_fpu_cp_req_valid),
    .io_fpu_cp_req_bits_cmd(core_io_fpu_cp_req_bits_cmd),
    .io_fpu_cp_req_bits_ldst(core_io_fpu_cp_req_bits_ldst),
    .io_fpu_cp_req_bits_wen(core_io_fpu_cp_req_bits_wen),
    .io_fpu_cp_req_bits_ren1(core_io_fpu_cp_req_bits_ren1),
    .io_fpu_cp_req_bits_ren2(core_io_fpu_cp_req_bits_ren2),
    .io_fpu_cp_req_bits_ren3(core_io_fpu_cp_req_bits_ren3),
    .io_fpu_cp_req_bits_swap12(core_io_fpu_cp_req_bits_swap12),
    .io_fpu_cp_req_bits_swap23(core_io_fpu_cp_req_bits_swap23),
    .io_fpu_cp_req_bits_single(core_io_fpu_cp_req_bits_single),
    .io_fpu_cp_req_bits_fromint(core_io_fpu_cp_req_bits_fromint),
    .io_fpu_cp_req_bits_toint(core_io_fpu_cp_req_bits_toint),
    .io_fpu_cp_req_bits_fastpipe(core_io_fpu_cp_req_bits_fastpipe),
    .io_fpu_cp_req_bits_fma(core_io_fpu_cp_req_bits_fma),
    .io_fpu_cp_req_bits_div(core_io_fpu_cp_req_bits_div),
    .io_fpu_cp_req_bits_sqrt(core_io_fpu_cp_req_bits_sqrt),
    .io_fpu_cp_req_bits_round(core_io_fpu_cp_req_bits_round),
    .io_fpu_cp_req_bits_wflags(core_io_fpu_cp_req_bits_wflags),
    .io_fpu_cp_req_bits_rm(core_io_fpu_cp_req_bits_rm),
    .io_fpu_cp_req_bits_typ(core_io_fpu_cp_req_bits_typ),
    .io_fpu_cp_req_bits_in1(core_io_fpu_cp_req_bits_in1),
    .io_fpu_cp_req_bits_in2(core_io_fpu_cp_req_bits_in2),
    .io_fpu_cp_req_bits_in3(core_io_fpu_cp_req_bits_in3),
    .io_fpu_cp_resp_ready(core_io_fpu_cp_resp_ready),
    .io_fpu_cp_resp_valid(core_io_fpu_cp_resp_valid),
    .io_fpu_cp_resp_bits_data(core_io_fpu_cp_resp_bits_data),
    .io_fpu_cp_resp_bits_exc(core_io_fpu_cp_resp_bits_exc),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(core_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(core_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(core_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(core_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(core_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(core_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(core_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(core_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(core_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(core_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(core_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(core_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(core_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(core_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(core_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(core_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(core_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(core_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(core_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(core_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(core_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(core_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(core_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(core_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(core_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(core_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(core_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(core_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(core_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(core_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(core_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(core_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(core_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(core_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(core_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(core_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(core_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(core_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(core_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(core_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(core_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(core_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(core_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(core_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(core_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(core_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(core_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(core_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(core_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(core_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(core_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(core_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(core_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(core_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(core_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(core_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(core_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(core_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(core_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(core_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(core_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(core_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(core_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(core_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(core_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(core_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(core_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(core_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(core_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(core_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(core_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(core_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(core_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(core_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(core_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(core_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(core_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(core_io_rocc_exception),
    .io_rocc_csr_waddr(core_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(core_io_rocc_csr_wdata),
    .io_rocc_csr_wen(core_io_rocc_csr_wen),
    .io_rocc_host_id(core_io_rocc_host_id)
  );
  
  //<CJ> RESET_VECTOR_ADDR
   defparam icache.RESET_VECTOR_ADDR = RESET_VECTOR_ADDR;
  
  CORERISCV_AXI4_FRONTEND icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_pc(icache_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(icache_io_cpu_req_bits_speculative),
    .io_cpu_resp_ready(icache_io_cpu_resp_ready),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(icache_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data_0(icache_io_cpu_resp_bits_data_0),
    .io_cpu_resp_bits_mask(icache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_if(icache_io_cpu_resp_bits_xcpt_if),
    .io_cpu_resp_bits_replay(icache_io_cpu_resp_bits_replay),
    .io_cpu_btb_resp_valid(icache_io_cpu_btb_resp_valid),
    .io_cpu_btb_resp_bits_taken(icache_io_cpu_btb_resp_bits_taken),
    .io_cpu_btb_resp_bits_mask(icache_io_cpu_btb_resp_bits_mask),
    .io_cpu_btb_resp_bits_bridx(icache_io_cpu_btb_resp_bits_bridx),
    .io_cpu_btb_resp_bits_target(icache_io_cpu_btb_resp_bits_target),
    .io_cpu_btb_resp_bits_entry(icache_io_cpu_btb_resp_bits_entry),
    .io_cpu_btb_resp_bits_bht_history(icache_io_cpu_btb_resp_bits_bht_history),
    .io_cpu_btb_resp_bits_bht_value(icache_io_cpu_btb_resp_bits_bht_value),
    .io_cpu_btb_update_valid(icache_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_valid(icache_io_cpu_btb_update_bits_prediction_valid),
    .io_cpu_btb_update_bits_prediction_bits_taken(icache_io_cpu_btb_update_bits_prediction_bits_taken),
    .io_cpu_btb_update_bits_prediction_bits_mask(icache_io_cpu_btb_update_bits_prediction_bits_mask),
    .io_cpu_btb_update_bits_prediction_bits_bridx(icache_io_cpu_btb_update_bits_prediction_bits_bridx),
    .io_cpu_btb_update_bits_prediction_bits_target(icache_io_cpu_btb_update_bits_prediction_bits_target),
    .io_cpu_btb_update_bits_prediction_bits_entry(icache_io_cpu_btb_update_bits_prediction_bits_entry),
    .io_cpu_btb_update_bits_prediction_bits_bht_history(icache_io_cpu_btb_update_bits_prediction_bits_bht_history),
    .io_cpu_btb_update_bits_prediction_bits_bht_value(icache_io_cpu_btb_update_bits_prediction_bits_bht_value),
    .io_cpu_btb_update_bits_pc(icache_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_target(icache_io_cpu_btb_update_bits_target),
    .io_cpu_btb_update_bits_taken(icache_io_cpu_btb_update_bits_taken),
    .io_cpu_btb_update_bits_isJump(icache_io_cpu_btb_update_bits_isJump),
    .io_cpu_btb_update_bits_isReturn(icache_io_cpu_btb_update_bits_isReturn),
    .io_cpu_btb_update_bits_br_pc(icache_io_cpu_btb_update_bits_br_pc),
    .io_cpu_bht_update_valid(icache_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_valid(icache_io_cpu_bht_update_bits_prediction_valid),
    .io_cpu_bht_update_bits_prediction_bits_taken(icache_io_cpu_bht_update_bits_prediction_bits_taken),
    .io_cpu_bht_update_bits_prediction_bits_mask(icache_io_cpu_bht_update_bits_prediction_bits_mask),
    .io_cpu_bht_update_bits_prediction_bits_bridx(icache_io_cpu_bht_update_bits_prediction_bits_bridx),
    .io_cpu_bht_update_bits_prediction_bits_target(icache_io_cpu_bht_update_bits_prediction_bits_target),
    .io_cpu_bht_update_bits_prediction_bits_entry(icache_io_cpu_bht_update_bits_prediction_bits_entry),
    .io_cpu_bht_update_bits_prediction_bits_bht_history(icache_io_cpu_bht_update_bits_prediction_bits_bht_history),
    .io_cpu_bht_update_bits_prediction_bits_bht_value(icache_io_cpu_bht_update_bits_prediction_bits_bht_value),
    .io_cpu_bht_update_bits_pc(icache_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_taken(icache_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(icache_io_cpu_bht_update_bits_mispredict),
    .io_cpu_ras_update_valid(icache_io_cpu_ras_update_valid),
    .io_cpu_ras_update_bits_isCall(icache_io_cpu_ras_update_bits_isCall),
    .io_cpu_ras_update_bits_isReturn(icache_io_cpu_ras_update_bits_isReturn),
    .io_cpu_ras_update_bits_returnAddr(icache_io_cpu_ras_update_bits_returnAddr),
    .io_cpu_ras_update_bits_prediction_valid(icache_io_cpu_ras_update_bits_prediction_valid),
    .io_cpu_ras_update_bits_prediction_bits_taken(icache_io_cpu_ras_update_bits_prediction_bits_taken),
    .io_cpu_ras_update_bits_prediction_bits_mask(icache_io_cpu_ras_update_bits_prediction_bits_mask),
    .io_cpu_ras_update_bits_prediction_bits_bridx(icache_io_cpu_ras_update_bits_prediction_bits_bridx),
    .io_cpu_ras_update_bits_prediction_bits_target(icache_io_cpu_ras_update_bits_prediction_bits_target),
    .io_cpu_ras_update_bits_prediction_bits_entry(icache_io_cpu_ras_update_bits_prediction_bits_entry),
    .io_cpu_ras_update_bits_prediction_bits_bht_history(icache_io_cpu_ras_update_bits_prediction_bits_bht_history),
    .io_cpu_ras_update_bits_prediction_bits_bht_value(icache_io_cpu_ras_update_bits_prediction_bits_bht_value),
    .io_cpu_flush_icache(icache_io_cpu_flush_icache),
    .io_cpu_flush_tlb(icache_io_cpu_flush_tlb),
    .io_cpu_npc(icache_io_cpu_npc),
    .io_ptw_req_ready(icache_io_ptw_req_ready),
    .io_ptw_req_valid(icache_io_ptw_req_valid),
    .io_ptw_req_bits_prv(icache_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(icache_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(icache_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(icache_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(icache_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(icache_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(icache_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(icache_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(icache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(icache_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(icache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(icache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(icache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(icache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(icache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(icache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(icache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(icache_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(icache_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(icache_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(icache_io_ptw_invalidate),
    .io_ptw_status_debug(icache_io_ptw_status_debug),
    .io_ptw_status_prv(icache_io_ptw_status_prv),
    .io_ptw_status_sd(icache_io_ptw_status_sd),
    .io_ptw_status_zero3(icache_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(icache_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(icache_io_ptw_status_zero2),
    .io_ptw_status_vm(icache_io_ptw_status_vm),
    .io_ptw_status_zero1(icache_io_ptw_status_zero1),
    .io_ptw_status_mxr(icache_io_ptw_status_mxr),
    .io_ptw_status_pum(icache_io_ptw_status_pum),
    .io_ptw_status_mprv(icache_io_ptw_status_mprv),
    .io_ptw_status_xs(icache_io_ptw_status_xs),
    .io_ptw_status_fs(icache_io_ptw_status_fs),
    .io_ptw_status_mpp(icache_io_ptw_status_mpp),
    .io_ptw_status_hpp(icache_io_ptw_status_hpp),
    .io_ptw_status_spp(icache_io_ptw_status_spp),
    .io_ptw_status_mpie(icache_io_ptw_status_mpie),
    .io_ptw_status_hpie(icache_io_ptw_status_hpie),
    .io_ptw_status_spie(icache_io_ptw_status_spie),
    .io_ptw_status_upie(icache_io_ptw_status_upie),
    .io_ptw_status_mie(icache_io_ptw_status_mie),
    .io_ptw_status_hie(icache_io_ptw_status_hie),
    .io_ptw_status_sie(icache_io_ptw_status_sie),
    .io_ptw_status_uie(icache_io_ptw_status_uie),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  CORERISCV_AXI4_D_CACHE DCache_1 (
    .clk(DCache_1_clk),
    .reset(DCache_1_reset),
    .io_cpu_req_ready(DCache_1_io_cpu_req_ready),
    .io_cpu_req_valid(DCache_1_io_cpu_req_valid),
    .io_cpu_req_bits_addr(DCache_1_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(DCache_1_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(DCache_1_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(DCache_1_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(DCache_1_io_cpu_req_bits_phys),
    .io_cpu_req_bits_data(DCache_1_io_cpu_req_bits_data),
    .io_cpu_s1_kill(DCache_1_io_cpu_s1_kill),
    .io_cpu_s1_data(DCache_1_io_cpu_s1_data),
    .io_cpu_s2_nack(DCache_1_io_cpu_s2_nack),
    .io_cpu_resp_valid(DCache_1_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(DCache_1_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(DCache_1_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(DCache_1_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_typ(DCache_1_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(DCache_1_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(DCache_1_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(DCache_1_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(DCache_1_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_store_data(DCache_1_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(DCache_1_io_cpu_replay_next),
    .io_cpu_xcpt_ma_ld(DCache_1_io_cpu_xcpt_ma_ld),
    .io_cpu_xcpt_ma_st(DCache_1_io_cpu_xcpt_ma_st),
    .io_cpu_xcpt_pf_ld(DCache_1_io_cpu_xcpt_pf_ld),
    .io_cpu_xcpt_pf_st(DCache_1_io_cpu_xcpt_pf_st),
    .io_cpu_invalidate_lr(DCache_1_io_cpu_invalidate_lr),
    .io_cpu_ordered(DCache_1_io_cpu_ordered),
    .io_ptw_req_ready(DCache_1_io_ptw_req_ready),
    .io_ptw_req_valid(DCache_1_io_ptw_req_valid),
    .io_ptw_req_bits_prv(DCache_1_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(DCache_1_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(DCache_1_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(DCache_1_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(DCache_1_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(DCache_1_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(DCache_1_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(DCache_1_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(DCache_1_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(DCache_1_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(DCache_1_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(DCache_1_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(DCache_1_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(DCache_1_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(DCache_1_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(DCache_1_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(DCache_1_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(DCache_1_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(DCache_1_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(DCache_1_io_ptw_invalidate),
    .io_ptw_status_debug(DCache_1_io_ptw_status_debug),
    .io_ptw_status_prv(DCache_1_io_ptw_status_prv),
    .io_ptw_status_sd(DCache_1_io_ptw_status_sd),
    .io_ptw_status_zero3(DCache_1_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(DCache_1_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(DCache_1_io_ptw_status_zero2),
    .io_ptw_status_vm(DCache_1_io_ptw_status_vm),
    .io_ptw_status_zero1(DCache_1_io_ptw_status_zero1),
    .io_ptw_status_mxr(DCache_1_io_ptw_status_mxr),
    .io_ptw_status_pum(DCache_1_io_ptw_status_pum),
    .io_ptw_status_mprv(DCache_1_io_ptw_status_mprv),
    .io_ptw_status_xs(DCache_1_io_ptw_status_xs),
    .io_ptw_status_fs(DCache_1_io_ptw_status_fs),
    .io_ptw_status_mpp(DCache_1_io_ptw_status_mpp),
    .io_ptw_status_hpp(DCache_1_io_ptw_status_hpp),
    .io_ptw_status_spp(DCache_1_io_ptw_status_spp),
    .io_ptw_status_mpie(DCache_1_io_ptw_status_mpie),
    .io_ptw_status_hpie(DCache_1_io_ptw_status_hpie),
    .io_ptw_status_spie(DCache_1_io_ptw_status_spie),
    .io_ptw_status_upie(DCache_1_io_ptw_status_upie),
    .io_ptw_status_mie(DCache_1_io_ptw_status_mie),
    .io_ptw_status_hie(DCache_1_io_ptw_status_hie),
    .io_ptw_status_sie(DCache_1_io_ptw_status_sie),
    .io_ptw_status_uie(DCache_1_io_ptw_status_uie),
    .io_mem_acquire_ready(DCache_1_io_mem_acquire_ready),
    .io_mem_acquire_valid(DCache_1_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(DCache_1_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(DCache_1_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(DCache_1_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(DCache_1_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(DCache_1_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(DCache_1_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(DCache_1_io_mem_acquire_bits_data),
    .io_mem_probe_ready(DCache_1_io_mem_probe_ready),
    .io_mem_probe_valid(DCache_1_io_mem_probe_valid),
    .io_mem_probe_bits_addr_block(DCache_1_io_mem_probe_bits_addr_block),
    .io_mem_probe_bits_p_type(DCache_1_io_mem_probe_bits_p_type),
    .io_mem_release_ready(DCache_1_io_mem_release_ready),
    .io_mem_release_valid(DCache_1_io_mem_release_valid),
    .io_mem_release_bits_addr_beat(DCache_1_io_mem_release_bits_addr_beat),
    .io_mem_release_bits_addr_block(DCache_1_io_mem_release_bits_addr_block),
    .io_mem_release_bits_client_xact_id(DCache_1_io_mem_release_bits_client_xact_id),
    .io_mem_release_bits_voluntary(DCache_1_io_mem_release_bits_voluntary),
    .io_mem_release_bits_r_type(DCache_1_io_mem_release_bits_r_type),
    .io_mem_release_bits_data(DCache_1_io_mem_release_bits_data),
    .io_mem_grant_ready(DCache_1_io_mem_grant_ready),
    .io_mem_grant_valid(DCache_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(DCache_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(DCache_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(DCache_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(DCache_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(DCache_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(DCache_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(DCache_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(DCache_1_io_mem_finish_ready),
    .io_mem_finish_valid(DCache_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(DCache_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(DCache_1_io_mem_finish_bits_manager_id)
  );
  CORERISCV_AXI4_CLIENT_UNCACHED_TILE_LINK_IO_ARBITER uncachedArb (
    .clk(uncachedArb_clk),
    .reset(uncachedArb_reset),
    .io_in_0_acquire_ready(uncachedArb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(uncachedArb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(uncachedArb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(uncachedArb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(uncachedArb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(uncachedArb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(uncachedArb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(uncachedArb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(uncachedArb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(uncachedArb_io_in_0_grant_ready),
    .io_in_0_grant_valid(uncachedArb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(uncachedArb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(uncachedArb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(uncachedArb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(uncachedArb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(uncachedArb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(uncachedArb_io_in_0_grant_bits_data),
    .io_out_acquire_ready(uncachedArb_io_out_acquire_ready),
    .io_out_acquire_valid(uncachedArb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(uncachedArb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(uncachedArb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(uncachedArb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(uncachedArb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(uncachedArb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(uncachedArb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(uncachedArb_io_out_acquire_bits_data),
    .io_out_grant_ready(uncachedArb_io_out_grant_ready),
    .io_out_grant_valid(uncachedArb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(uncachedArb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(uncachedArb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(uncachedArb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(uncachedArb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(uncachedArb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(uncachedArb_io_out_grant_bits_data)
  );
  CORERISCV_AXI4_HELLA_CACHE_ARBITER dcArb (
    .clk(dcArb_clk),
    .reset(dcArb_reset),
    .io_requestor_0_req_ready(dcArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_data(dcArb_io_requestor_0_req_bits_data),
    .io_requestor_0_s1_kill(dcArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data(dcArb_io_requestor_0_s1_data),
    .io_requestor_0_s2_nack(dcArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(dcArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(dcArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(dcArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_typ(dcArb_io_requestor_0_resp_bits_typ),
    .io_requestor_0_resp_bits_data(dcArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_replay(dcArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(dcArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(dcArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_store_data(dcArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(dcArb_io_requestor_0_replay_next),
    .io_requestor_0_xcpt_ma_ld(dcArb_io_requestor_0_xcpt_ma_ld),
    .io_requestor_0_xcpt_ma_st(dcArb_io_requestor_0_xcpt_ma_st),
    .io_requestor_0_xcpt_pf_ld(dcArb_io_requestor_0_xcpt_pf_ld),
    .io_requestor_0_xcpt_pf_st(dcArb_io_requestor_0_xcpt_pf_st),
    .io_requestor_0_invalidate_lr(dcArb_io_requestor_0_invalidate_lr),
    .io_requestor_0_ordered(dcArb_io_requestor_0_ordered),
    .io_mem_req_ready(dcArb_io_mem_req_ready),
    .io_mem_req_valid(dcArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcArb_io_mem_req_bits_phys),
    .io_mem_req_bits_data(dcArb_io_mem_req_bits_data),
    .io_mem_s1_kill(dcArb_io_mem_s1_kill),
    .io_mem_s1_data(dcArb_io_mem_s1_data),
    .io_mem_s2_nack(dcArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(dcArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(dcArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(dcArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(dcArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(dcArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(dcArb_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(dcArb_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(dcArb_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(dcArb_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(dcArb_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(dcArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcArb_io_mem_ordered)
  );
  assign io_cached_0_acquire_valid = DCache_1_io_mem_acquire_valid;
  assign io_cached_0_acquire_bits_addr_block = DCache_1_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_bits_client_xact_id = DCache_1_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_beat = DCache_1_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_is_builtin_type = DCache_1_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_a_type = DCache_1_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_union = DCache_1_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_data = DCache_1_io_mem_acquire_bits_data;
  assign io_cached_0_probe_ready = DCache_1_io_mem_probe_ready;
  assign io_cached_0_release_valid = DCache_1_io_mem_release_valid;
  assign io_cached_0_release_bits_addr_beat = DCache_1_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_bits_addr_block = DCache_1_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_client_xact_id = DCache_1_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_voluntary = DCache_1_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = DCache_1_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_data = DCache_1_io_mem_release_bits_data;
  assign io_cached_0_grant_ready = DCache_1_io_mem_grant_ready;
  assign io_cached_0_finish_valid = DCache_1_io_mem_finish_valid;
  assign io_cached_0_finish_bits_manager_xact_id = DCache_1_io_mem_finish_bits_manager_xact_id;
  assign io_cached_0_finish_bits_manager_id = DCache_1_io_mem_finish_bits_manager_id;
  assign io_uncached_0_acquire_valid = uncachedArb_io_out_acquire_valid;
  assign io_uncached_0_acquire_bits_addr_block = uncachedArb_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_bits_client_xact_id = uncachedArb_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_beat = uncachedArb_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_is_builtin_type = uncachedArb_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_a_type = uncachedArb_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_union = uncachedArb_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_data = uncachedArb_io_out_acquire_bits_data;
  assign io_uncached_0_grant_ready = uncachedArb_io_out_grant_ready;
  assign core_clk = clk;
  assign core_reset = reset;
  assign core_io_prci_reset = io_prci_reset;
  assign core_io_prci_id = io_prci_id;
  assign core_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign core_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign core_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign core_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign core_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign core_io_imem_resp_valid = icache_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_pc = icache_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data_0 = icache_io_cpu_resp_bits_data_0;
  assign core_io_imem_resp_bits_mask = icache_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_if = icache_io_cpu_resp_bits_xcpt_if;
  assign core_io_imem_resp_bits_replay = icache_io_cpu_resp_bits_replay;
  assign core_io_imem_btb_resp_valid = icache_io_cpu_btb_resp_valid;
  assign core_io_imem_btb_resp_bits_taken = icache_io_cpu_btb_resp_bits_taken;
  assign core_io_imem_btb_resp_bits_mask = icache_io_cpu_btb_resp_bits_mask;
  assign core_io_imem_btb_resp_bits_bridx = icache_io_cpu_btb_resp_bits_bridx;
  assign core_io_imem_btb_resp_bits_target = icache_io_cpu_btb_resp_bits_target;
  assign core_io_imem_btb_resp_bits_entry = icache_io_cpu_btb_resp_bits_entry;
  assign core_io_imem_btb_resp_bits_bht_history = icache_io_cpu_btb_resp_bits_bht_history;
  assign core_io_imem_btb_resp_bits_bht_value = icache_io_cpu_btb_resp_bits_bht_value;
  assign core_io_imem_npc = icache_io_cpu_npc;
  assign core_io_dmem_req_ready = dcArb_io_requestor_0_req_ready;
  assign core_io_dmem_s2_nack = dcArb_io_requestor_0_s2_nack;
  assign core_io_dmem_resp_valid = dcArb_io_requestor_0_resp_valid;
  assign core_io_dmem_resp_bits_addr = dcArb_io_requestor_0_resp_bits_addr;
  assign core_io_dmem_resp_bits_tag = dcArb_io_requestor_0_resp_bits_tag;
  assign core_io_dmem_resp_bits_cmd = dcArb_io_requestor_0_resp_bits_cmd;
  assign core_io_dmem_resp_bits_typ = dcArb_io_requestor_0_resp_bits_typ;
  assign core_io_dmem_resp_bits_data = dcArb_io_requestor_0_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcArb_io_requestor_0_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcArb_io_requestor_0_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcArb_io_requestor_0_resp_bits_data_word_bypass;
  assign core_io_dmem_resp_bits_store_data = dcArb_io_requestor_0_resp_bits_store_data;
  assign core_io_dmem_replay_next = dcArb_io_requestor_0_replay_next;
  assign core_io_dmem_xcpt_ma_ld = dcArb_io_requestor_0_xcpt_ma_ld;
  assign core_io_dmem_xcpt_ma_st = dcArb_io_requestor_0_xcpt_ma_st;
  assign core_io_dmem_xcpt_pf_ld = dcArb_io_requestor_0_xcpt_pf_ld;
  assign core_io_dmem_xcpt_pf_st = dcArb_io_requestor_0_xcpt_pf_st;
  assign core_io_dmem_ordered = dcArb_io_requestor_0_ordered;
  assign core_io_fpu_fcsr_flags_valid = GEN_0;
  assign core_io_fpu_fcsr_flags_bits = GEN_1;
  assign core_io_fpu_store_data = GEN_2;
  assign core_io_fpu_toint_data = GEN_3;
  assign core_io_fpu_fcsr_rdy = GEN_4;
  assign core_io_fpu_nack_mem = GEN_5;
  assign core_io_fpu_illegal_rm = GEN_6;
  assign core_io_fpu_dec_cmd = GEN_7;
  assign core_io_fpu_dec_ldst = GEN_8;
  assign core_io_fpu_dec_wen = GEN_9;
  assign core_io_fpu_dec_ren1 = GEN_10;
  assign core_io_fpu_dec_ren2 = GEN_11;
  assign core_io_fpu_dec_ren3 = GEN_12;
  assign core_io_fpu_dec_swap12 = GEN_13;
  assign core_io_fpu_dec_swap23 = GEN_14;
  assign core_io_fpu_dec_single = GEN_15;
  assign core_io_fpu_dec_fromint = GEN_16;
  assign core_io_fpu_dec_toint = GEN_17;
  assign core_io_fpu_dec_fastpipe = GEN_18;
  assign core_io_fpu_dec_fma = GEN_19;
  assign core_io_fpu_dec_div = GEN_20;
  assign core_io_fpu_dec_sqrt = GEN_21;
  assign core_io_fpu_dec_round = GEN_22;
  assign core_io_fpu_dec_wflags = GEN_23;
  assign core_io_fpu_sboard_set = GEN_24;
  assign core_io_fpu_sboard_clr = GEN_25;
  assign core_io_fpu_sboard_clra = GEN_26;
  assign core_io_fpu_cp_req_ready = GEN_27;
  assign core_io_fpu_cp_resp_valid = GEN_28;
  assign core_io_fpu_cp_resp_bits_data = GEN_29;
  assign core_io_fpu_cp_resp_bits_exc = GEN_30;
  assign core_io_rocc_cmd_ready = GEN_31;
  assign core_io_rocc_resp_valid = GEN_32;
  assign core_io_rocc_resp_bits_rd = GEN_33;
  assign core_io_rocc_resp_bits_data = GEN_34;
  assign core_io_rocc_mem_req_valid = GEN_35;
  assign core_io_rocc_mem_req_bits_addr = GEN_36;
  assign core_io_rocc_mem_req_bits_tag = GEN_37;
  assign core_io_rocc_mem_req_bits_cmd = GEN_38;
  assign core_io_rocc_mem_req_bits_typ = GEN_39;
  assign core_io_rocc_mem_req_bits_phys = GEN_40;
  assign core_io_rocc_mem_req_bits_data = GEN_41;
  assign core_io_rocc_mem_s1_kill = GEN_42;
  assign core_io_rocc_mem_s1_data = GEN_43;
  assign core_io_rocc_mem_invalidate_lr = GEN_44;
  assign core_io_rocc_busy = GEN_45;
  assign core_io_rocc_interrupt = GEN_46;
  assign core_io_rocc_autl_acquire_valid = GEN_47;
  assign core_io_rocc_autl_acquire_bits_addr_block = GEN_48;
  assign core_io_rocc_autl_acquire_bits_client_xact_id = GEN_49;
  assign core_io_rocc_autl_acquire_bits_addr_beat = GEN_50;
  assign core_io_rocc_autl_acquire_bits_is_builtin_type = GEN_51;
  assign core_io_rocc_autl_acquire_bits_a_type = GEN_52;
  assign core_io_rocc_autl_acquire_bits_union = GEN_53;
  assign core_io_rocc_autl_acquire_bits_data = GEN_54;
  assign core_io_rocc_autl_grant_ready = GEN_55;
  assign core_io_rocc_fpu_req_valid = GEN_56;
  assign core_io_rocc_fpu_req_bits_cmd = GEN_57;
  assign core_io_rocc_fpu_req_bits_ldst = GEN_58;
  assign core_io_rocc_fpu_req_bits_wen = GEN_59;
  assign core_io_rocc_fpu_req_bits_ren1 = GEN_60;
  assign core_io_rocc_fpu_req_bits_ren2 = GEN_61;
  assign core_io_rocc_fpu_req_bits_ren3 = GEN_62;
  assign core_io_rocc_fpu_req_bits_swap12 = GEN_63;
  assign core_io_rocc_fpu_req_bits_swap23 = GEN_64;
  assign core_io_rocc_fpu_req_bits_single = GEN_65;
  assign core_io_rocc_fpu_req_bits_fromint = GEN_66;
  assign core_io_rocc_fpu_req_bits_toint = GEN_67;
  assign core_io_rocc_fpu_req_bits_fastpipe = GEN_68;
  assign core_io_rocc_fpu_req_bits_fma = GEN_69;
  assign core_io_rocc_fpu_req_bits_div = GEN_70;
  assign core_io_rocc_fpu_req_bits_sqrt = GEN_71;
  assign core_io_rocc_fpu_req_bits_round = GEN_72;
  assign core_io_rocc_fpu_req_bits_wflags = GEN_73;
  assign core_io_rocc_fpu_req_bits_rm = GEN_74;
  assign core_io_rocc_fpu_req_bits_typ = GEN_75;
  assign core_io_rocc_fpu_req_bits_in1 = GEN_76;
  assign core_io_rocc_fpu_req_bits_in2 = GEN_77;
  assign core_io_rocc_fpu_req_bits_in3 = GEN_78;
  assign core_io_rocc_fpu_resp_ready = GEN_79;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_cpu_req_valid = core_io_imem_req_valid;
  assign icache_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign icache_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
  assign icache_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign icache_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
  assign icache_io_cpu_btb_update_bits_prediction_valid = core_io_imem_btb_update_bits_prediction_valid;
  assign icache_io_cpu_btb_update_bits_prediction_bits_taken = core_io_imem_btb_update_bits_prediction_bits_taken;
  assign icache_io_cpu_btb_update_bits_prediction_bits_mask = core_io_imem_btb_update_bits_prediction_bits_mask;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bridx = core_io_imem_btb_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_btb_update_bits_prediction_bits_target = core_io_imem_btb_update_bits_prediction_bits_target;
  assign icache_io_cpu_btb_update_bits_prediction_bits_entry = core_io_imem_btb_update_bits_prediction_bits_entry;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_history = core_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_value = core_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
  assign icache_io_cpu_btb_update_bits_target = core_io_imem_btb_update_bits_target;
  assign icache_io_cpu_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
  assign icache_io_cpu_btb_update_bits_isJump = core_io_imem_btb_update_bits_isJump;
  assign icache_io_cpu_btb_update_bits_isReturn = core_io_imem_btb_update_bits_isReturn;
  assign icache_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
  assign icache_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
  assign icache_io_cpu_bht_update_bits_prediction_valid = core_io_imem_bht_update_bits_prediction_valid;
  assign icache_io_cpu_bht_update_bits_prediction_bits_taken = core_io_imem_bht_update_bits_prediction_bits_taken;
  assign icache_io_cpu_bht_update_bits_prediction_bits_mask = core_io_imem_bht_update_bits_prediction_bits_mask;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bridx = core_io_imem_bht_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_bht_update_bits_prediction_bits_target = core_io_imem_bht_update_bits_prediction_bits_target;
  assign icache_io_cpu_bht_update_bits_prediction_bits_entry = core_io_imem_bht_update_bits_prediction_bits_entry;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_history = core_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_value = core_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
  assign icache_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
  assign icache_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
  assign icache_io_cpu_ras_update_valid = core_io_imem_ras_update_valid;
  assign icache_io_cpu_ras_update_bits_isCall = core_io_imem_ras_update_bits_isCall;
  assign icache_io_cpu_ras_update_bits_isReturn = core_io_imem_ras_update_bits_isReturn;
  assign icache_io_cpu_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
  assign icache_io_cpu_ras_update_bits_prediction_valid = core_io_imem_ras_update_bits_prediction_valid;
  assign icache_io_cpu_ras_update_bits_prediction_bits_taken = core_io_imem_ras_update_bits_prediction_bits_taken;
  assign icache_io_cpu_ras_update_bits_prediction_bits_mask = core_io_imem_ras_update_bits_prediction_bits_mask;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bridx = core_io_imem_ras_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_ras_update_bits_prediction_bits_target = core_io_imem_ras_update_bits_prediction_bits_target;
  assign icache_io_cpu_ras_update_bits_prediction_bits_entry = core_io_imem_ras_update_bits_prediction_bits_entry;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_history = core_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_value = core_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign icache_io_cpu_flush_tlb = core_io_imem_flush_tlb;
  assign icache_io_ptw_req_ready = GEN_80;
  assign icache_io_ptw_resp_valid = GEN_81;
  assign icache_io_ptw_resp_bits_pte_reserved_for_hardware = GEN_82;
  assign icache_io_ptw_resp_bits_pte_ppn = GEN_83;
  assign icache_io_ptw_resp_bits_pte_reserved_for_software = GEN_84;
  assign icache_io_ptw_resp_bits_pte_d = GEN_85;
  assign icache_io_ptw_resp_bits_pte_a = GEN_86;
  assign icache_io_ptw_resp_bits_pte_g = GEN_87;
  assign icache_io_ptw_resp_bits_pte_u = GEN_88;
  assign icache_io_ptw_resp_bits_pte_x = GEN_89;
  assign icache_io_ptw_resp_bits_pte_w = GEN_90;
  assign icache_io_ptw_resp_bits_pte_r = GEN_91;
  assign icache_io_ptw_resp_bits_pte_v = GEN_92;
  assign icache_io_ptw_ptbr_asid = GEN_93;
  assign icache_io_ptw_ptbr_ppn = GEN_94;
  assign icache_io_ptw_invalidate = GEN_95;
  assign icache_io_ptw_status_debug = GEN_96;
  assign icache_io_ptw_status_prv = GEN_97;
  assign icache_io_ptw_status_sd = GEN_98;
  assign icache_io_ptw_status_zero3 = GEN_99;
  assign icache_io_ptw_status_sd_rv32 = GEN_100;
  assign icache_io_ptw_status_zero2 = GEN_101;
  assign icache_io_ptw_status_vm = GEN_102;
  assign icache_io_ptw_status_zero1 = GEN_103;
  assign icache_io_ptw_status_mxr = GEN_104;
  assign icache_io_ptw_status_pum = GEN_105;
  assign icache_io_ptw_status_mprv = GEN_106;
  assign icache_io_ptw_status_xs = GEN_107;
  assign icache_io_ptw_status_fs = GEN_108;
  assign icache_io_ptw_status_mpp = GEN_109;
  assign icache_io_ptw_status_hpp = GEN_110;
  assign icache_io_ptw_status_spp = GEN_111;
  assign icache_io_ptw_status_mpie = GEN_112;
  assign icache_io_ptw_status_hpie = GEN_113;
  assign icache_io_ptw_status_spie = GEN_114;
  assign icache_io_ptw_status_upie = GEN_115;
  assign icache_io_ptw_status_mie = GEN_116;
  assign icache_io_ptw_status_hie = GEN_117;
  assign icache_io_ptw_status_sie = GEN_118;
  assign icache_io_ptw_status_uie = GEN_119;
  assign icache_io_mem_acquire_ready = uncachedArb_io_in_0_acquire_ready;
  assign icache_io_mem_grant_valid = uncachedArb_io_in_0_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = uncachedArb_io_in_0_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = uncachedArb_io_in_0_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = uncachedArb_io_in_0_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = uncachedArb_io_in_0_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = uncachedArb_io_in_0_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = uncachedArb_io_in_0_grant_bits_data;
  assign DCache_1_clk = clk;
  assign DCache_1_reset = reset;
  assign DCache_1_io_cpu_req_valid = dcArb_io_mem_req_valid;
  assign DCache_1_io_cpu_req_bits_addr = dcArb_io_mem_req_bits_addr;
  assign DCache_1_io_cpu_req_bits_tag = dcArb_io_mem_req_bits_tag;
  assign DCache_1_io_cpu_req_bits_cmd = dcArb_io_mem_req_bits_cmd;
  assign DCache_1_io_cpu_req_bits_typ = dcArb_io_mem_req_bits_typ;
  assign DCache_1_io_cpu_req_bits_phys = dcArb_io_mem_req_bits_phys;
  assign DCache_1_io_cpu_req_bits_data = dcArb_io_mem_req_bits_data;
  assign DCache_1_io_cpu_s1_kill = dcArb_io_mem_s1_kill;
  assign DCache_1_io_cpu_s1_data = dcArb_io_mem_s1_data;
  assign DCache_1_io_cpu_invalidate_lr = dcArb_io_mem_invalidate_lr;
  assign DCache_1_io_ptw_req_ready = GEN_120;
  assign DCache_1_io_ptw_resp_valid = GEN_121;
  assign DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware = GEN_122;
  assign DCache_1_io_ptw_resp_bits_pte_ppn = GEN_123;
  assign DCache_1_io_ptw_resp_bits_pte_reserved_for_software = GEN_124;
  assign DCache_1_io_ptw_resp_bits_pte_d = GEN_125;
  assign DCache_1_io_ptw_resp_bits_pte_a = GEN_126;
  assign DCache_1_io_ptw_resp_bits_pte_g = GEN_127;
  assign DCache_1_io_ptw_resp_bits_pte_u = GEN_128;
  assign DCache_1_io_ptw_resp_bits_pte_x = GEN_129;
  assign DCache_1_io_ptw_resp_bits_pte_w = GEN_130;
  assign DCache_1_io_ptw_resp_bits_pte_r = GEN_131;
  assign DCache_1_io_ptw_resp_bits_pte_v = GEN_132;
  assign DCache_1_io_ptw_ptbr_asid = GEN_133;
  assign DCache_1_io_ptw_ptbr_ppn = GEN_134;
  assign DCache_1_io_ptw_invalidate = GEN_135;
  assign DCache_1_io_ptw_status_debug = GEN_136;
  assign DCache_1_io_ptw_status_prv = GEN_137;
  assign DCache_1_io_ptw_status_sd = GEN_138;
  assign DCache_1_io_ptw_status_zero3 = GEN_139;
  assign DCache_1_io_ptw_status_sd_rv32 = GEN_140;
  assign DCache_1_io_ptw_status_zero2 = GEN_141;
  assign DCache_1_io_ptw_status_vm = GEN_142;
  assign DCache_1_io_ptw_status_zero1 = GEN_143;
  assign DCache_1_io_ptw_status_mxr = GEN_144;
  assign DCache_1_io_ptw_status_pum = GEN_145;
  assign DCache_1_io_ptw_status_mprv = GEN_146;
  assign DCache_1_io_ptw_status_xs = GEN_147;
  assign DCache_1_io_ptw_status_fs = GEN_148;
  assign DCache_1_io_ptw_status_mpp = GEN_149;
  assign DCache_1_io_ptw_status_hpp = GEN_150;
  assign DCache_1_io_ptw_status_spp = GEN_151;
  assign DCache_1_io_ptw_status_mpie = GEN_152;
  assign DCache_1_io_ptw_status_hpie = GEN_153;
  assign DCache_1_io_ptw_status_spie = GEN_154;
  assign DCache_1_io_ptw_status_upie = GEN_155;
  assign DCache_1_io_ptw_status_mie = GEN_156;
  assign DCache_1_io_ptw_status_hie = GEN_157;
  assign DCache_1_io_ptw_status_sie = GEN_158;
  assign DCache_1_io_ptw_status_uie = GEN_159;
  assign DCache_1_io_mem_acquire_ready = io_cached_0_acquire_ready;
  assign DCache_1_io_mem_probe_valid = io_cached_0_probe_valid;
  assign DCache_1_io_mem_probe_bits_addr_block = io_cached_0_probe_bits_addr_block;
  assign DCache_1_io_mem_probe_bits_p_type = io_cached_0_probe_bits_p_type;
  assign DCache_1_io_mem_release_ready = io_cached_0_release_ready;
  assign DCache_1_io_mem_grant_valid = io_cached_0_grant_valid;
  assign DCache_1_io_mem_grant_bits_addr_beat = io_cached_0_grant_bits_addr_beat;
  assign DCache_1_io_mem_grant_bits_client_xact_id = io_cached_0_grant_bits_client_xact_id;
  assign DCache_1_io_mem_grant_bits_manager_xact_id = io_cached_0_grant_bits_manager_xact_id;
  assign DCache_1_io_mem_grant_bits_is_builtin_type = io_cached_0_grant_bits_is_builtin_type;
  assign DCache_1_io_mem_grant_bits_g_type = io_cached_0_grant_bits_g_type;
  assign DCache_1_io_mem_grant_bits_data = io_cached_0_grant_bits_data;
  assign DCache_1_io_mem_grant_bits_manager_id = io_cached_0_grant_bits_manager_id;
  assign DCache_1_io_mem_finish_ready = io_cached_0_finish_ready;
  assign uncachedArb_clk = clk;
  assign uncachedArb_reset = reset;
  assign uncachedArb_io_in_0_acquire_valid = icache_io_mem_acquire_valid;
  assign uncachedArb_io_in_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign uncachedArb_io_in_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign uncachedArb_io_in_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign uncachedArb_io_in_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign uncachedArb_io_in_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign uncachedArb_io_in_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign uncachedArb_io_in_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign uncachedArb_io_in_0_grant_ready = icache_io_mem_grant_ready;
  assign uncachedArb_io_out_acquire_ready = io_uncached_0_acquire_ready;
  assign uncachedArb_io_out_grant_valid = io_uncached_0_grant_valid;
  assign uncachedArb_io_out_grant_bits_addr_beat = io_uncached_0_grant_bits_addr_beat;
  assign uncachedArb_io_out_grant_bits_client_xact_id = io_uncached_0_grant_bits_client_xact_id;
  assign uncachedArb_io_out_grant_bits_manager_xact_id = io_uncached_0_grant_bits_manager_xact_id;
  assign uncachedArb_io_out_grant_bits_is_builtin_type = io_uncached_0_grant_bits_is_builtin_type;
  assign uncachedArb_io_out_grant_bits_g_type = io_uncached_0_grant_bits_g_type;
  assign uncachedArb_io_out_grant_bits_data = io_uncached_0_grant_bits_data;
  assign dcArb_clk = clk;
  assign dcArb_reset = reset;
  assign dcArb_io_requestor_0_req_valid = core_io_dmem_req_valid;
  assign dcArb_io_requestor_0_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcArb_io_requestor_0_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcArb_io_requestor_0_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcArb_io_requestor_0_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcArb_io_requestor_0_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcArb_io_requestor_0_req_bits_data = core_io_dmem_req_bits_data;
  assign dcArb_io_requestor_0_s1_kill = core_io_dmem_s1_kill;
  assign dcArb_io_requestor_0_s1_data = core_io_dmem_s1_data;
  assign dcArb_io_requestor_0_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcArb_io_mem_req_ready = DCache_1_io_cpu_req_ready;
  assign dcArb_io_mem_s2_nack = DCache_1_io_cpu_s2_nack;
  assign dcArb_io_mem_resp_valid = DCache_1_io_cpu_resp_valid;
  assign dcArb_io_mem_resp_bits_addr = DCache_1_io_cpu_resp_bits_addr;
  assign dcArb_io_mem_resp_bits_tag = DCache_1_io_cpu_resp_bits_tag;
  assign dcArb_io_mem_resp_bits_cmd = DCache_1_io_cpu_resp_bits_cmd;
  assign dcArb_io_mem_resp_bits_typ = DCache_1_io_cpu_resp_bits_typ;
  assign dcArb_io_mem_resp_bits_data = DCache_1_io_cpu_resp_bits_data;
  assign dcArb_io_mem_resp_bits_replay = DCache_1_io_cpu_resp_bits_replay;
  assign dcArb_io_mem_resp_bits_has_data = DCache_1_io_cpu_resp_bits_has_data;
  assign dcArb_io_mem_resp_bits_data_word_bypass = DCache_1_io_cpu_resp_bits_data_word_bypass;
  assign dcArb_io_mem_resp_bits_store_data = DCache_1_io_cpu_resp_bits_store_data;
  assign dcArb_io_mem_replay_next = DCache_1_io_cpu_replay_next;
  assign dcArb_io_mem_xcpt_ma_ld = DCache_1_io_cpu_xcpt_ma_ld;
  assign dcArb_io_mem_xcpt_ma_st = DCache_1_io_cpu_xcpt_ma_st;
  assign dcArb_io_mem_xcpt_pf_ld = DCache_1_io_cpu_xcpt_pf_ld;
  assign dcArb_io_mem_xcpt_pf_st = DCache_1_io_cpu_xcpt_pf_st;
  assign dcArb_io_mem_ordered = DCache_1_io_cpu_ordered;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_160 = {1{$random}};
  GEN_0 = GEN_160[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_161 = {1{$random}};
  GEN_1 = GEN_161[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_162 = {2{$random}};
  GEN_2 = GEN_162[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_163 = {1{$random}};
  GEN_3 = GEN_163[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_164 = {1{$random}};
  GEN_4 = GEN_164[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_165 = {1{$random}};
  GEN_5 = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_166 = {1{$random}};
  GEN_6 = GEN_166[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_167 = {1{$random}};
  GEN_7 = GEN_167[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_168 = {1{$random}};
  GEN_8 = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_169 = {1{$random}};
  GEN_9 = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_170 = {1{$random}};
  GEN_10 = GEN_170[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_171 = {1{$random}};
  GEN_11 = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_172 = {1{$random}};
  GEN_12 = GEN_172[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_173 = {1{$random}};
  GEN_13 = GEN_173[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_174 = {1{$random}};
  GEN_14 = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_175 = {1{$random}};
  GEN_15 = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_176 = {1{$random}};
  GEN_16 = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_177 = {1{$random}};
  GEN_17 = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_178 = {1{$random}};
  GEN_18 = GEN_178[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_179 = {1{$random}};
  GEN_19 = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_180 = {1{$random}};
  GEN_20 = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_181 = {1{$random}};
  GEN_21 = GEN_181[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_182 = {1{$random}};
  GEN_22 = GEN_182[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_183 = {1{$random}};
  GEN_23 = GEN_183[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_184 = {1{$random}};
  GEN_24 = GEN_184[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_185 = {1{$random}};
  GEN_25 = GEN_185[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_186 = {1{$random}};
  GEN_26 = GEN_186[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_187 = {1{$random}};
  GEN_27 = GEN_187[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_188 = {1{$random}};
  GEN_28 = GEN_188[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_189 = {3{$random}};
  GEN_29 = GEN_189[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_190 = {1{$random}};
  GEN_30 = GEN_190[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_191 = {1{$random}};
  GEN_31 = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_192 = {1{$random}};
  GEN_32 = GEN_192[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_193 = {1{$random}};
  GEN_33 = GEN_193[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_194 = {1{$random}};
  GEN_34 = GEN_194[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_195 = {1{$random}};
  GEN_35 = GEN_195[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_196 = {1{$random}};
  GEN_36 = GEN_196[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_197 = {1{$random}};
  GEN_37 = GEN_197[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_198 = {1{$random}};
  GEN_38 = GEN_198[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_199 = {1{$random}};
  GEN_39 = GEN_199[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_200 = {1{$random}};
  GEN_40 = GEN_200[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_201 = {1{$random}};
  GEN_41 = GEN_201[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_202 = {1{$random}};
  GEN_42 = GEN_202[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_203 = {1{$random}};
  GEN_43 = GEN_203[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_204 = {1{$random}};
  GEN_44 = GEN_204[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_205 = {1{$random}};
  GEN_45 = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_206 = {1{$random}};
  GEN_46 = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_207 = {1{$random}};
  GEN_47 = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_208 = {1{$random}};
  GEN_48 = GEN_208[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_209 = {1{$random}};
  GEN_49 = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_210 = {1{$random}};
  GEN_50 = GEN_210[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_211 = {1{$random}};
  GEN_51 = GEN_211[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_212 = {1{$random}};
  GEN_52 = GEN_212[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_213 = {1{$random}};
  GEN_53 = GEN_213[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_214 = {2{$random}};
  GEN_54 = GEN_214[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_215 = {1{$random}};
  GEN_55 = GEN_215[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_216 = {1{$random}};
  GEN_56 = GEN_216[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_217 = {1{$random}};
  GEN_57 = GEN_217[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_218 = {1{$random}};
  GEN_58 = GEN_218[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_219 = {1{$random}};
  GEN_59 = GEN_219[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_220 = {1{$random}};
  GEN_60 = GEN_220[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_221 = {1{$random}};
  GEN_61 = GEN_221[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_222 = {1{$random}};
  GEN_62 = GEN_222[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_223 = {1{$random}};
  GEN_63 = GEN_223[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_224 = {1{$random}};
  GEN_64 = GEN_224[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_225 = {1{$random}};
  GEN_65 = GEN_225[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_226 = {1{$random}};
  GEN_66 = GEN_226[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_227 = {1{$random}};
  GEN_67 = GEN_227[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_228 = {1{$random}};
  GEN_68 = GEN_228[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_229 = {1{$random}};
  GEN_69 = GEN_229[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_230 = {1{$random}};
  GEN_70 = GEN_230[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_231 = {1{$random}};
  GEN_71 = GEN_231[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_232 = {1{$random}};
  GEN_72 = GEN_232[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_233 = {1{$random}};
  GEN_73 = GEN_233[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_234 = {1{$random}};
  GEN_74 = GEN_234[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_235 = {1{$random}};
  GEN_75 = GEN_235[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_236 = {3{$random}};
  GEN_76 = GEN_236[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_237 = {3{$random}};
  GEN_77 = GEN_237[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_238 = {3{$random}};
  GEN_78 = GEN_238[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_239 = {1{$random}};
  GEN_79 = GEN_239[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_240 = {1{$random}};
  GEN_80 = GEN_240[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_241 = {1{$random}};
  GEN_81 = GEN_241[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_242 = {1{$random}};
  GEN_82 = GEN_242[15:0];
  `endif
  `ifdef RANDOMIZE
  GEN_243 = {2{$random}};
  GEN_83 = GEN_243[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_244 = {1{$random}};
  GEN_84 = GEN_244[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_245 = {1{$random}};
  GEN_85 = GEN_245[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_246 = {1{$random}};
  GEN_86 = GEN_246[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_247 = {1{$random}};
  GEN_87 = GEN_247[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_248 = {1{$random}};
  GEN_88 = GEN_248[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_249 = {1{$random}};
  GEN_89 = GEN_249[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_250 = {1{$random}};
  GEN_90 = GEN_250[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_251 = {1{$random}};
  GEN_91 = GEN_251[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_252 = {1{$random}};
  GEN_92 = GEN_252[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_253 = {1{$random}};
  GEN_93 = GEN_253[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_254 = {1{$random}};
  GEN_94 = GEN_254[21:0];
  `endif
  `ifdef RANDOMIZE
  GEN_255 = {1{$random}};
  GEN_95 = GEN_255[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_256 = {1{$random}};
  GEN_96 = GEN_256[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_257 = {1{$random}};
  GEN_97 = GEN_257[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_258 = {1{$random}};
  GEN_98 = GEN_258[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_259 = {1{$random}};
  GEN_99 = GEN_259[30:0];
  `endif
  `ifdef RANDOMIZE
  GEN_260 = {1{$random}};
  GEN_100 = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_261 = {1{$random}};
  GEN_101 = GEN_261[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_262 = {1{$random}};
  GEN_102 = GEN_262[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_263 = {1{$random}};
  GEN_103 = GEN_263[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_264 = {1{$random}};
  GEN_104 = GEN_264[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_265 = {1{$random}};
  GEN_105 = GEN_265[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_266 = {1{$random}};
  GEN_106 = GEN_266[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_267 = {1{$random}};
  GEN_107 = GEN_267[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_268 = {1{$random}};
  GEN_108 = GEN_268[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_269 = {1{$random}};
  GEN_109 = GEN_269[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_270 = {1{$random}};
  GEN_110 = GEN_270[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_271 = {1{$random}};
  GEN_111 = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_272 = {1{$random}};
  GEN_112 = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_273 = {1{$random}};
  GEN_113 = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_274 = {1{$random}};
  GEN_114 = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_275 = {1{$random}};
  GEN_115 = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_276 = {1{$random}};
  GEN_116 = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_277 = {1{$random}};
  GEN_117 = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_278 = {1{$random}};
  GEN_118 = GEN_278[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_279 = {1{$random}};
  GEN_119 = GEN_279[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_280 = {1{$random}};
  GEN_120 = GEN_280[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_281 = {1{$random}};
  GEN_121 = GEN_281[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_282 = {1{$random}};
  GEN_122 = GEN_282[15:0];
  `endif
  `ifdef RANDOMIZE
  GEN_283 = {2{$random}};
  GEN_123 = GEN_283[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_284 = {1{$random}};
  GEN_124 = GEN_284[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_285 = {1{$random}};
  GEN_125 = GEN_285[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_286 = {1{$random}};
  GEN_126 = GEN_286[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_287 = {1{$random}};
  GEN_127 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_288 = {1{$random}};
  GEN_128 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_289 = {1{$random}};
  GEN_129 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_290 = {1{$random}};
  GEN_130 = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_291 = {1{$random}};
  GEN_131 = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_292 = {1{$random}};
  GEN_132 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_293 = {1{$random}};
  GEN_133 = GEN_293[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_294 = {1{$random}};
  GEN_134 = GEN_294[21:0];
  `endif
  `ifdef RANDOMIZE
  GEN_295 = {1{$random}};
  GEN_135 = GEN_295[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_296 = {1{$random}};
  GEN_136 = GEN_296[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_297 = {1{$random}};
  GEN_137 = GEN_297[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_298 = {1{$random}};
  GEN_138 = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_299 = {1{$random}};
  GEN_139 = GEN_299[30:0];
  `endif
  `ifdef RANDOMIZE
  GEN_300 = {1{$random}};
  GEN_140 = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_301 = {1{$random}};
  GEN_141 = GEN_301[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_302 = {1{$random}};
  GEN_142 = GEN_302[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_303 = {1{$random}};
  GEN_143 = GEN_303[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_304 = {1{$random}};
  GEN_144 = GEN_304[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_305 = {1{$random}};
  GEN_145 = GEN_305[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_306 = {1{$random}};
  GEN_146 = GEN_306[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_307 = {1{$random}};
  GEN_147 = GEN_307[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_308 = {1{$random}};
  GEN_148 = GEN_308[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_309 = {1{$random}};
  GEN_149 = GEN_309[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_310 = {1{$random}};
  GEN_150 = GEN_310[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_311 = {1{$random}};
  GEN_151 = GEN_311[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_312 = {1{$random}};
  GEN_152 = GEN_312[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_313 = {1{$random}};
  GEN_153 = GEN_313[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_314 = {1{$random}};
  GEN_154 = GEN_314[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_315 = {1{$random}};
  GEN_155 = GEN_315[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_316 = {1{$random}};
  GEN_156 = GEN_316[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_317 = {1{$random}};
  GEN_157 = GEN_317[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_318 = {1{$random}};
  GEN_158 = GEN_318[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_319 = {1{$random}};
  GEN_159 = GEN_319[0:0];
  `endif
  end
`endif
endmodule
